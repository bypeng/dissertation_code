module ntt8192_163841 ( clk, rst, start, input_fg, addr, din, dout, valid );

  localparam Q0 = 163841;

  // STATE
  localparam ST_IDLE   = 0;
  localparam ST_NTT    = 1;
  localparam ST_PMUL   = 2;
  localparam ST_RELOAD = 3;
  localparam ST_INTT   = 4;
  localparam ST_CRT    = 5;  // not applied for single prime scheme
  localparam ST_REDUCE = 6;
  localparam ST_FINISH = 7;

  input                      clk;
  input                      rst;
  input                      start;
  input                      input_fg;
  input             [13 : 0] addr;
  input signed      [17 : 0] din;
  output reg signed [17 : 0] dout;
  output reg                 valid;

  // BRAM
  reg            wr_en   [0 : 1];
  reg   [13 : 0] wr_addr [0 : 1];
  reg   [13 : 0] rd_addr [0 : 1];
  reg   [17 : 0] wr_din  [0 : 1];
  wire  [17 : 0] rd_dout [0 : 1];
  wire  [17 : 0] wr_dout [0 : 1];

  // addr_gen
  wire         bank_index_rd [0 : 1];
  wire         bank_index_wr [0 : 1];
  wire [12: 0] data_index_rd [0 : 1];
  wire [12: 0] data_index_wr [0 : 1];
  reg  bank_index_wr_0_shift_1, bank_index_wr_0_shift_2;
  reg  fg_shift_1, fg_shift_2, fg_shift_3;

  // w_addr_gen
  reg  [12 : 0] stage_bit;
  wire [12 : 0] w_addr;

  // bfu
  reg                  ntt_state; 
  reg  signed [17: 0] in_a  ;
  reg  signed [17: 0] in_b  ;
  reg  signed [17: 0] in_w  ;
  wire signed [35: 0] bw    ;
  wire signed [17: 0] out_a ;
  wire signed [17: 0] out_b ;

  // state, stage, counter
  reg  [2 : 0] state, next_state;
  reg  [4 : 0] stage, stage_wr;
  wire [4 : 0] stage_rdM, stage_wrM;
  reg  [14 : 0] ctr;
  reg  [14 : 0] ctr_shift_7, ctr_shift_8, ctr_shift_9, ctr_shift_1, ctr_shift_2;
  reg          ctr_MSB_masked;
  reg          poly_select;
  reg          ctr_msb_shift_1;
  wire         ctr_half_end, ctr_full_end, ctr_shift_7_end, stage_rd_end, stage_rd_2, stage_wr_end, ntt_end, point_proc_end, reduce_end;

  // w_array
  reg         [13: 0] w_addr_in;
  wire signed [17: 0] w_dout ;

  // misc
  reg          bank_index_rd_shift_1, bank_index_rd_shift_2;
  reg [13: 0] wr_ctr [0 : 1];
  reg [17: 0] din_shift_1, din_shift_2, din_shift_3;
  reg [13: 0] w_addr_in_shift_1;

  // BRAM instances
  bram_18_14_P bank_0
  (clk, wr_en[0], wr_addr[0], rd_addr[0], wr_din[0], wr_dout[0], rd_dout[0]);
  bram_18_14_P bank_1
  (clk, wr_en[1], wr_addr[1], rd_addr[1], wr_din[1], wr_dout[1], rd_dout[1]);

  // Read/Write Address Generator
  addr_gen addr_rd_0 (clk, stage_rdM, {ctr_MSB_masked, ctr[12:0]}, bank_index_rd[0], data_index_rd[0]);
  addr_gen addr_rd_1 (clk, stage_rdM, {1'b1, ctr[12:0]}, bank_index_rd[1], data_index_rd[1]);
  addr_gen addr_wr_0 (clk, stage_wrM, {wr_ctr[0]}, bank_index_wr[0], data_index_wr[0]);
  addr_gen addr_wr_1 (clk, stage_wrM, {wr_ctr[1]}, bank_index_wr[1], data_index_wr[1]);

  // Omega Address Generator
  w_addr_gen w_addr_gen_0 (clk, stage_bit, ctr[12:0], w_addr);

  // Butterfly Unit  , each with a corresponding omega array
  bfu_163841 bfu_inst (clk, ntt_state, in_a, in_b, in_w, bw, out_a, out_b);
  w_163841 rom_w_inst (clk, w_addr_in_shift_1, w_dout);

  assign ctr_half_end         = (ctr[12:0] == 8191) ? 1 : 0;
  assign ctr_full_end         = (ctr[13:0] == 16383) ? 1 : 0;
  assign stage_rd_end         = (stage == 14) ? 1 : 0;
  assign stage_rd_2           = (stage == 2) ? 1 : 0;
  assign ntt_end         = (stage_rd_end && ctr[12 : 0] == 10) ? 1 : 0;
  assign crt_end         = (stage_rd_2 && ctr[12 : 0] == 10) ? 1 : 0;
  assign point_proc_end   = (ctr == 16394) ? 1 : 0;
  assign reload_end      = (stage != 0 && ctr[12:0] == 4) ? 1 : 0;
  assign reduce_end      = (ctr == 16388);

  // crt
  // fg_shift
  always @ ( posedge clk ) begin
    fg_shift_1 <= input_fg;
    fg_shift_2 <= fg_shift_1;
    fg_shift_3 <= fg_shift_2;
  end
  // dout
  always @ ( posedge clk ) begin
    if (state == ST_FINISH) begin
      if (bank_index_wr_0_shift_2) begin
        dout <= wr_dout[1][17:0];
      end else begin
        dout <= wr_dout[0][17:0];
      end
    end else begin
      dout <= 'sd0;
    end
  end

  // bank_index_wr_0_shift_1
  always @ ( posedge clk ) begin
    bank_index_wr_0_shift_1 <= bank_index_wr[0];
    bank_index_wr_0_shift_2 <= bank_index_wr_0_shift_1;
  end

  // poly_select
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        poly_select <= ~poly_select;
      end else begin
        poly_select <= poly_select;
      end    
    end else if (state == ST_RELOAD) begin
      poly_select <= 1;
    end else begin
      poly_select <= 0;
    end
  end

  // w_addr_in_shift_1
  always @ ( posedge clk ) begin
    w_addr_in_shift_1 <= w_addr_in;
  end

  // din_shift
  always @ ( posedge clk ) begin
    din_shift_1 <= din;
    din_shift_2 <= din_shift_1;
    din_shift_3 <= din_shift_2;
  end

  // rd_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_rd[0]) begin
        rd_addr[0][12:0] <= data_index_rd[1];
        rd_addr[1][12:0] <= data_index_rd[0];
      end else begin
        rd_addr[0][12:0] <= data_index_rd[0];
        rd_addr[1][12:0] <= data_index_rd[1];
      end
    end else begin
      rd_addr[0][12:0] <= data_index_rd[0];
      rd_addr[1][12:0] <= data_index_rd[0];
    end

    if (state == ST_NTT)  begin
      rd_addr[0][13] <= poly_select;
      rd_addr[1][13] <= poly_select;
    end else if (state == ST_PMUL) begin
      rd_addr[0][13] <=  bank_index_rd[0];
      rd_addr[1][13] <= ~bank_index_rd[0];
    end else if (state == ST_RELOAD) begin
      rd_addr[0][13] <= 0;
      rd_addr[1][13] <= 0;
    end else begin
      rd_addr[0][13] <= 1;
      rd_addr[1][13] <= 1;
    end
  end

  // wr_en
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 1;
      end
    end else if (state == ST_IDLE) begin
      if (fg_shift_3 ^ bank_index_wr[0]) begin
        wr_en[0] <= 0;
        wr_en[1] <= 1;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 0;
      end
    end else if (state == ST_PMUL) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_REDUCE) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_CRT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else if (state == ST_RELOAD) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else begin
      wr_en[0] <= 0;
      wr_en[1] <= 0;
    end
  end

  // wr_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_addr[0][12:0] <= data_index_wr[1];
        wr_addr[1][12:0] <= data_index_wr[0];
      end else begin
        wr_addr[0][12:0] <= data_index_wr[0];
        wr_addr[1][12:0] <= data_index_wr[1];
      end
    end else begin
      wr_addr[0][12:0] <= data_index_wr[0];
      wr_addr[1][12:0] <= data_index_wr[0];
    end  

    if (state == ST_IDLE) begin
      wr_addr[0][13] <= fg_shift_3;
      wr_addr[1][13] <= fg_shift_3;
    end else if(state == ST_NTT || state == ST_INTT) begin
      wr_addr[0][13] <= poly_select;
      wr_addr[1][13] <= poly_select;
    end else if (state == ST_PMUL || state == ST_REDUCE || state == ST_FINISH) begin
      wr_addr[0][13] <= 0;
      wr_addr[1][13] <= 0;
    end else begin
      wr_addr[0][13] <= 1;
      wr_addr[1][13] <= 1;
    end     
  end

  // wr_din
  always @ ( posedge clk ) begin
    if (state == ST_IDLE) begin
      wr_din[0][17:0] <= { din_shift_3 };
      wr_din[1][17:0] <= { din_shift_3 };
    end else if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_din[0][17:0] <= out_b;
        wr_din[1][17:0] <= out_a;
      end else begin
        wr_din[0][17:0] <= out_a;
        wr_din[1][17:0] <= out_b;
      end
    end else if (state == ST_RELOAD) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end
    end else if (state == ST_REDUCE) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end
    end else begin
      wr_din[0][17:0] <= out_a;
      wr_din[1][17:0] <= out_a;
    end
  end

  // bank_index_rd_shift
  always @ ( posedge clk ) begin
    bank_index_rd_shift_1 <= bank_index_rd[0];
    bank_index_rd_shift_2 <= bank_index_rd_shift_1;
  end

  // ntt_state
  always @ ( posedge clk ) begin
    if (state == ST_INTT) begin
      ntt_state <= 1;
    end else begin
      ntt_state <= 0;
    end
  end

  // in_a, in_b
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else if (state == ST_CRT) begin
      if (bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else begin // ST_PMUL
      in_b <= $signed(rd_dout[1]);
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_a <= $signed(rd_dout[1]);
      end else begin
        in_a <= $signed(rd_dout[0]);
      end
    end else begin // ST_PMUL, ST_CRT
      in_a <= 'sd0;
    end
  end

  // w_addr_in, in_w
  always @ ( posedge clk ) begin
    if (state == ST_NTT) begin
      w_addr_in <= {1'b0, w_addr};
    end else begin
      w_addr_in <= 16384 - w_addr;
    end

    if (state == ST_PMUL) begin
        in_w <= rd_dout[0];
    end else begin
      in_w <= w_dout;
    end
  end

  // wr_ctr
  always @ ( posedge clk ) begin
    if (state == ST_IDLE || state == ST_FINISH) begin
      wr_ctr[0] <= addr[13:0];
    end else if (state == ST_RELOAD || state == ST_REDUCE) begin
      wr_ctr[0] <= {ctr_shift_1[0], ctr_shift_1[1], ctr_shift_1[2], ctr_shift_1[3], ctr_shift_1[4], ctr_shift_1[5], ctr_shift_1[6], ctr_shift_1[7], ctr_shift_1[8], ctr_shift_1[9], ctr_shift_1[10], ctr_shift_1[11], ctr_shift_1[12], ctr_shift_1[13]};
    end else if (state == ST_NTT || state == ST_INTT) begin
      wr_ctr[0] <= {1'b0, ctr_shift_7[12:0]};
    end else begin
      wr_ctr[0] <= ctr_shift_7[13:0];
    end

    wr_ctr[1] <= {1'b1, ctr_shift_7[12:0]};
  end

  // ctr_MSB_masked
  always @ (*) begin
    if (state == ST_NTT || state == ST_INTT) begin
      ctr_MSB_masked = 0;
    end else begin
      ctr_MSB_masked = ctr[13];
    end
  end

  // ctr, ctr_shifts
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_PMUL) begin
      if (point_proc_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_CRT) begin
      if (crt_end || ctr_full_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_REDUCE) begin
      if (reduce_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else begin
      ctr <= 0;
    end

    //change ctr_shift_7 <= ctr - 5;
    ctr_shift_7 <= ctr - 7;
    ctr_shift_8 <= ctr_shift_7;
    ctr_shift_9 <= ctr_shift_8;
    ctr_shift_1 <= ctr;
    ctr_shift_2 <= ctr_shift_1;
  end

  // stage, stage_wr
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage <= 0;
      end else if (ctr_half_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else begin
      stage <= 0;
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[12:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[13:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_9[13:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else begin
      stage_wr <= 0;
    end        
  end
  assign stage_rdM = (state == ST_NTT || state == ST_INTT) ? stage : 0;
  assign stage_wrM = (state == ST_NTT || state == ST_INTT) ? stage_wr : 0;

  // stage_bit
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_bit <= 0;
      end else if (ctr_half_end) begin
        stage_bit[0] <= 1'b1;
        stage_bit[12 : 1] <= stage_bit[11 : 0];
      end else begin
        stage_bit <= stage_bit;
      end
    end else begin
      stage_bit <= 'b0;
    end
  end

  // valid
  always @ (*) begin
      if (state == ST_FINISH) begin
          valid = 1;
      end else begin
          valid = 0;
      end
  end

  // state
  always @ ( posedge clk ) begin
    if(rst) begin
            state <= 0;
        end else begin
            state <= next_state;
        end
  end

  always @(*) begin
    case(state)
    ST_IDLE: begin
      if(start)
        next_state = ST_NTT;
      else
        next_state = ST_IDLE;
    end
    ST_NTT: begin
      if(ntt_end && poly_select == 1)
        next_state = ST_PMUL;
      else
        next_state = ST_NTT;
    end
    ST_PMUL: begin
      if (point_proc_end)
        next_state = ST_RELOAD;
      else
        next_state = ST_PMUL;
    end
    ST_RELOAD: begin
      if (reload_end) begin
        next_state = ST_INTT;
      end else begin
        next_state = ST_RELOAD;
      end
    end
    ST_INTT: begin
      if(ntt_end)
        next_state = ST_REDUCE;
      else
        next_state = ST_INTT;
      end
    ST_REDUCE: begin
      if(reduce_end)
        next_state = ST_FINISH;
      else
        next_state = ST_REDUCE;
    end
    ST_FINISH: begin
      if(!start)
        next_state = ST_FINISH;
      else
        next_state = ST_IDLE;
    end
    default: next_state = ST_IDLE;
    endcase
  end

endmodule

module w_addr_gen ( clk, stage_bit, ctr, w_addr );

  input              clk;
  input      [12: 0] stage_bit;
  input      [12: 0] ctr;
  output reg [12: 0] w_addr;

  wire [12: 0] w;

  assign w[ 0] = (stage_bit[ 0]) ? ctr[ 0] : 0;
  assign w[ 1] = (stage_bit[ 1]) ? ctr[ 1] : 0;
  assign w[ 2] = (stage_bit[ 2]) ? ctr[ 2] : 0;
  assign w[ 3] = (stage_bit[ 3]) ? ctr[ 3] : 0;
  assign w[ 4] = (stage_bit[ 4]) ? ctr[ 4] : 0;
  assign w[ 5] = (stage_bit[ 5]) ? ctr[ 5] : 0;
  assign w[ 6] = (stage_bit[ 6]) ? ctr[ 6] : 0;
  assign w[ 7] = (stage_bit[ 7]) ? ctr[ 7] : 0;
  assign w[ 8] = (stage_bit[ 8]) ? ctr[ 8] : 0;
  assign w[ 9] = (stage_bit[ 9]) ? ctr[ 9] : 0;
  assign w[10] = (stage_bit[10]) ? ctr[10] : 0;
  assign w[11] = (stage_bit[11]) ? ctr[11] : 0;
  assign w[12] = (stage_bit[12]) ? ctr[12] : 0;

  always @ ( posedge clk ) begin
    w_addr <= {w[0], w[1], w[2], w[3], w[4], w[5], w[6], w[7], w[8], w[9], w[10], w[11], w[12]};
  end

endmodule

module addr_gen ( clk, stage, ctr, bank_index, data_index );

  input              clk;
  input      [3 : 0] stage;
  input      [13: 0] ctr;
  output reg         bank_index;
  output reg [12: 0] data_index;

  wire       [13: 0] bs_out;

  barrel_shifter bs ( clk, ctr, stage, bs_out );

    always @( posedge clk ) begin
        bank_index <= ^bs_out;
    end

    always @( posedge clk ) begin
        data_index <= bs_out[13:1];
    end

endmodule

module barrel_shifter ( clk, in, shift, out );

  input              clk;
  input      [13: 0] in;
  input      [3 : 0] shift;
  output reg [13: 0] out;

  reg        [13: 0] in_s [0:4];

  always @ (*) begin
    in_s[0] = in;
  end

  always @ (*) begin
    if(shift[0]) begin
      in_s[1] = { in_s[0][0], in_s[0][13:1] };
    end else begin
      in_s[1] = in_s[0];
    end
  end

  always @ (*) begin
    if(shift[1]) begin
      in_s[2] = { in_s[1][1:0], in_s[1][13:2] };
    end else begin
      in_s[2] = in_s[1];
    end
  end

  always @ (*) begin
    if(shift[2]) begin
      in_s[3] = { in_s[2][3:0], in_s[2][13:4] };
    end else begin
      in_s[3] = in_s[2];
    end
  end

  always @ (*) begin
    if(shift[3]) begin
      in_s[4] = { in_s[3][7:0], in_s[3][13:8] };
    end else begin
      in_s[4] = in_s[3];
    end
  end

  always @ ( posedge clk ) begin
    out <= in_s[4];
  end

endmodule

module bfu_163841 ( clk, state, in_a, in_b, w, bw, out_a, out_b );

  input                      clk;
  input                      state;
  input      signed [17 : 0] in_a;
  input      signed [17 : 0] in_b;
  input      signed [17 : 0] w;
  output reg signed [34 : 0] bw;
  output reg signed [17 : 0] out_a;
  output reg signed [17 : 0] out_b;

  wire signed       [17 : 0] mod_bw;
  reg signed        [18 : 0] a, b;
  reg signed        [17 : 0] in_a_s1, in_a_s2, in_a_s3, in_a_s4, in_a_s5;

  reg signed        [34 : 0] bwQ_0, bwQ_1, bwQ_2;
  wire signed       [18 : 0] a_add_q, a_sub_q, b_add_q, b_sub_q;

  modmul163841s mod163841s_inst ( clk, 1'b0, bw, mod_bw );

  assign a_add_q = a + 'sd163841;
  assign a_sub_q = a - 'sd163841;
  assign b_add_q = b + 'sd163841;
  assign b_sub_q = b - 'sd163841;

  always @(posedge clk ) begin
    in_a_s1 <= in_a;
    in_a_s2 <= in_a_s1;
    in_a_s3 <= in_a_s2;
    in_a_s4 <= in_a_s3;
    in_a_s5 <= in_a_s4;
  end

  always @ ( posedge clk ) begin
    bw <= in_b * w;
  end

  always @ ( posedge clk ) begin
    a <= in_a_s4 + mod_bw;
    b <= in_a_s4 - mod_bw;

    if (state == 0) begin
      if (a > 'sd81920) begin
        out_a <= a_sub_q;
      end else if (a < -'sd81920) begin
        out_a <= a_add_q;
      end else begin
        out_a <= a;
      end
    end else begin
      if (a[0] == 0) begin
        out_a <= a[18:1];
      end else if (a[18] == 0) begin // a > 0
        out_a <= a_sub_q[18:1];
      end else begin                 // a < 0
        out_a <= a_add_q[18:1];
      end
    end

    if (state == 0) begin
      if (b > 'sd81920) begin
        out_b <= b_sub_q;
      end else if (b < -'sd81920) begin
        out_b <= b_add_q;
      end else begin
        out_b <= b;
      end
    end else begin
      if (b[0] == 0) begin
        out_b <= b[18:1];
      end else if (b[18] == 0) begin // b > 0
        out_b <= b_sub_q[18:1];
      end else begin                 // b < 0
        out_b <= b_add_q[18:1];
      end
    end
  end

endmodule

module w_163841 ( clk, addr, dout );

  input                       clk;
  input             [13 : 0]  addr;
  output signed     [17 : 0]  dout;

  wire signed       [17 : 0]  dout_p;
  wire signed       [17 : 0]  dout_n;
  reg               [13 : 0]  addr_reg;

  (* rom_style = "block" *) reg signed [17:0] data [0:8191];

  assign dout_p = data[addr_reg[12:0]];
  assign dout_n = -dout_p;
  assign dout   = addr_reg[13] ? dout_n : dout_p;

  always @ ( posedge clk ) begin
    addr_reg <= addr;
  end

  initial begin
    data[   0] =  'sd1;
    data[   1] =  'sd5;
    data[   2] =  'sd25;
    data[   3] =  'sd125;
    data[   4] =  'sd625;
    data[   5] =  'sd3125;
    data[   6] =  'sd15625;
    data[   7] =  'sd78125;
    data[   8] =  'sd62943;
    data[   9] = -'sd12967;
    data[  10] = -'sd64835;
    data[  11] =  'sd3507;
    data[  12] =  'sd17535;
    data[  13] = -'sd76166;
    data[  14] = -'sd53148;
    data[  15] =  'sd61942;
    data[  16] = -'sd17972;
    data[  17] =  'sd73981;
    data[  18] =  'sd42223;
    data[  19] =  'sd47274;
    data[  20] =  'sd72529;
    data[  21] =  'sd34963;
    data[  22] =  'sd10974;
    data[  23] =  'sd54870;
    data[  24] = -'sd53332;
    data[  25] =  'sd61022;
    data[  26] = -'sd22572;
    data[  27] =  'sd50981;
    data[  28] = -'sd72777;
    data[  29] = -'sd36203;
    data[  30] = -'sd17174;
    data[  31] =  'sd77971;
    data[  32] =  'sd62173;
    data[  33] = -'sd16817;
    data[  34] =  'sd79756;
    data[  35] =  'sd71098;
    data[  36] =  'sd27808;
    data[  37] = -'sd24801;
    data[  38] =  'sd39836;
    data[  39] =  'sd35339;
    data[  40] =  'sd12854;
    data[  41] =  'sd64270;
    data[  42] = -'sd6332;
    data[  43] = -'sd31660;
    data[  44] =  'sd5541;
    data[  45] =  'sd27705;
    data[  46] = -'sd25316;
    data[  47] =  'sd37261;
    data[  48] =  'sd22464;
    data[  49] = -'sd51521;
    data[  50] =  'sd70077;
    data[  51] =  'sd22703;
    data[  52] = -'sd50326;
    data[  53] =  'sd76052;
    data[  54] =  'sd52578;
    data[  55] = -'sd64792;
    data[  56] =  'sd3722;
    data[  57] =  'sd18610;
    data[  58] = -'sd70791;
    data[  59] = -'sd26273;
    data[  60] =  'sd32476;
    data[  61] = -'sd1461;
    data[  62] = -'sd7305;
    data[  63] = -'sd36525;
    data[  64] = -'sd18784;
    data[  65] =  'sd69921;
    data[  66] =  'sd21923;
    data[  67] = -'sd54226;
    data[  68] =  'sd56552;
    data[  69] = -'sd44922;
    data[  70] = -'sd60769;
    data[  71] =  'sd23837;
    data[  72] = -'sd44656;
    data[  73] = -'sd59439;
    data[  74] =  'sd30487;
    data[  75] = -'sd11406;
    data[  76] = -'sd57030;
    data[  77] =  'sd42532;
    data[  78] =  'sd48819;
    data[  79] =  'sd80254;
    data[  80] =  'sd73588;
    data[  81] =  'sd40258;
    data[  82] =  'sd37449;
    data[  83] =  'sd23404;
    data[  84] = -'sd46821;
    data[  85] = -'sd70264;
    data[  86] = -'sd23638;
    data[  87] =  'sd45651;
    data[  88] =  'sd64414;
    data[  89] = -'sd5612;
    data[  90] = -'sd28060;
    data[  91] =  'sd23541;
    data[  92] = -'sd46136;
    data[  93] = -'sd66839;
    data[  94] = -'sd6513;
    data[  95] = -'sd32565;
    data[  96] =  'sd1016;
    data[  97] =  'sd5080;
    data[  98] =  'sd25400;
    data[  99] = -'sd36841;
    data[ 100] = -'sd20364;
    data[ 101] =  'sd62021;
    data[ 102] = -'sd17577;
    data[ 103] =  'sd75956;
    data[ 104] =  'sd52098;
    data[ 105] = -'sd67192;
    data[ 106] = -'sd8278;
    data[ 107] = -'sd41390;
    data[ 108] = -'sd43109;
    data[ 109] = -'sd51704;
    data[ 110] =  'sd69162;
    data[ 111] =  'sd18128;
    data[ 112] = -'sd73201;
    data[ 113] = -'sd38323;
    data[ 114] = -'sd27774;
    data[ 115] =  'sd24971;
    data[ 116] = -'sd38986;
    data[ 117] = -'sd31089;
    data[ 118] =  'sd8396;
    data[ 119] =  'sd41980;
    data[ 120] =  'sd46059;
    data[ 121] =  'sd66454;
    data[ 122] =  'sd4588;
    data[ 123] =  'sd22940;
    data[ 124] = -'sd49141;
    data[ 125] = -'sd81864;
    data[ 126] = -'sd81638;
    data[ 127] = -'sd80508;
    data[ 128] = -'sd74858;
    data[ 129] = -'sd46608;
    data[ 130] = -'sd69199;
    data[ 131] = -'sd18313;
    data[ 132] =  'sd72276;
    data[ 133] =  'sd33698;
    data[ 134] =  'sd4649;
    data[ 135] =  'sd23245;
    data[ 136] = -'sd47616;
    data[ 137] = -'sd74239;
    data[ 138] = -'sd43513;
    data[ 139] = -'sd53724;
    data[ 140] =  'sd59062;
    data[ 141] = -'sd32372;
    data[ 142] =  'sd1981;
    data[ 143] =  'sd9905;
    data[ 144] =  'sd49525;
    data[ 145] = -'sd80057;
    data[ 146] = -'sd72603;
    data[ 147] = -'sd35333;
    data[ 148] = -'sd12824;
    data[ 149] = -'sd64120;
    data[ 150] =  'sd7082;
    data[ 151] =  'sd35410;
    data[ 152] =  'sd13209;
    data[ 153] =  'sd66045;
    data[ 154] =  'sd2543;
    data[ 155] =  'sd12715;
    data[ 156] =  'sd63575;
    data[ 157] = -'sd9807;
    data[ 158] = -'sd49035;
    data[ 159] = -'sd81334;
    data[ 160] = -'sd78988;
    data[ 161] = -'sd67258;
    data[ 162] = -'sd8608;
    data[ 163] = -'sd43040;
    data[ 164] = -'sd51359;
    data[ 165] =  'sd70887;
    data[ 166] =  'sd26753;
    data[ 167] = -'sd30076;
    data[ 168] =  'sd13461;
    data[ 169] =  'sd67305;
    data[ 170] =  'sd8843;
    data[ 171] =  'sd44215;
    data[ 172] =  'sd57234;
    data[ 173] = -'sd41512;
    data[ 174] = -'sd43719;
    data[ 175] = -'sd54754;
    data[ 176] =  'sd53912;
    data[ 177] = -'sd58122;
    data[ 178] =  'sd37072;
    data[ 179] =  'sd21519;
    data[ 180] = -'sd56246;
    data[ 181] =  'sd46452;
    data[ 182] =  'sd68419;
    data[ 183] =  'sd14413;
    data[ 184] =  'sd72065;
    data[ 185] =  'sd32643;
    data[ 186] = -'sd626;
    data[ 187] = -'sd3130;
    data[ 188] = -'sd15650;
    data[ 189] = -'sd78250;
    data[ 190] = -'sd63568;
    data[ 191] =  'sd9842;
    data[ 192] =  'sd49210;
    data[ 193] = -'sd81632;
    data[ 194] = -'sd80478;
    data[ 195] = -'sd74708;
    data[ 196] = -'sd45858;
    data[ 197] = -'sd65449;
    data[ 198] =  'sd437;
    data[ 199] =  'sd2185;
    data[ 200] =  'sd10925;
    data[ 201] =  'sd54625;
    data[ 202] = -'sd54557;
    data[ 203] =  'sd54897;
    data[ 204] = -'sd53197;
    data[ 205] =  'sd61697;
    data[ 206] = -'sd19197;
    data[ 207] =  'sd67856;
    data[ 208] =  'sd11598;
    data[ 209] =  'sd57990;
    data[ 210] = -'sd37732;
    data[ 211] = -'sd24819;
    data[ 212] =  'sd39746;
    data[ 213] =  'sd34889;
    data[ 214] =  'sd10604;
    data[ 215] =  'sd53020;
    data[ 216] = -'sd62582;
    data[ 217] =  'sd14772;
    data[ 218] =  'sd73860;
    data[ 219] =  'sd41618;
    data[ 220] =  'sd44249;
    data[ 221] =  'sd57404;
    data[ 222] = -'sd40662;
    data[ 223] = -'sd39469;
    data[ 224] = -'sd33504;
    data[ 225] = -'sd3679;
    data[ 226] = -'sd18395;
    data[ 227] =  'sd71866;
    data[ 228] =  'sd31648;
    data[ 229] = -'sd5601;
    data[ 230] = -'sd28005;
    data[ 231] =  'sd23816;
    data[ 232] = -'sd44761;
    data[ 233] = -'sd59964;
    data[ 234] =  'sd27862;
    data[ 235] = -'sd24531;
    data[ 236] =  'sd41186;
    data[ 237] =  'sd42089;
    data[ 238] =  'sd46604;
    data[ 239] =  'sd69179;
    data[ 240] =  'sd18213;
    data[ 241] = -'sd72776;
    data[ 242] = -'sd36198;
    data[ 243] = -'sd17149;
    data[ 244] =  'sd78096;
    data[ 245] =  'sd62798;
    data[ 246] = -'sd13692;
    data[ 247] = -'sd68460;
    data[ 248] = -'sd14618;
    data[ 249] = -'sd73090;
    data[ 250] = -'sd37768;
    data[ 251] = -'sd24999;
    data[ 252] =  'sd38846;
    data[ 253] =  'sd30389;
    data[ 254] = -'sd11896;
    data[ 255] = -'sd59480;
    data[ 256] =  'sd30282;
    data[ 257] = -'sd12431;
    data[ 258] = -'sd62155;
    data[ 259] =  'sd16907;
    data[ 260] = -'sd79306;
    data[ 261] = -'sd68848;
    data[ 262] = -'sd16558;
    data[ 263] =  'sd81051;
    data[ 264] =  'sd77573;
    data[ 265] =  'sd60183;
    data[ 266] = -'sd26767;
    data[ 267] =  'sd30006;
    data[ 268] = -'sd13811;
    data[ 269] = -'sd69055;
    data[ 270] = -'sd17593;
    data[ 271] =  'sd75876;
    data[ 272] =  'sd51698;
    data[ 273] = -'sd69192;
    data[ 274] = -'sd18278;
    data[ 275] =  'sd72451;
    data[ 276] =  'sd34573;
    data[ 277] =  'sd9024;
    data[ 278] =  'sd45120;
    data[ 279] =  'sd61759;
    data[ 280] = -'sd18887;
    data[ 281] =  'sd69406;
    data[ 282] =  'sd19348;
    data[ 283] = -'sd67101;
    data[ 284] = -'sd7823;
    data[ 285] = -'sd39115;
    data[ 286] = -'sd31734;
    data[ 287] =  'sd5171;
    data[ 288] =  'sd25855;
    data[ 289] = -'sd34566;
    data[ 290] = -'sd8989;
    data[ 291] = -'sd44945;
    data[ 292] = -'sd60884;
    data[ 293] =  'sd23262;
    data[ 294] = -'sd47531;
    data[ 295] = -'sd73814;
    data[ 296] = -'sd41388;
    data[ 297] = -'sd43099;
    data[ 298] = -'sd51654;
    data[ 299] =  'sd69412;
    data[ 300] =  'sd19378;
    data[ 301] = -'sd66951;
    data[ 302] = -'sd7073;
    data[ 303] = -'sd35365;
    data[ 304] = -'sd12984;
    data[ 305] = -'sd64920;
    data[ 306] =  'sd3082;
    data[ 307] =  'sd15410;
    data[ 308] =  'sd77050;
    data[ 309] =  'sd57568;
    data[ 310] = -'sd39842;
    data[ 311] = -'sd35369;
    data[ 312] = -'sd13004;
    data[ 313] = -'sd65020;
    data[ 314] =  'sd2582;
    data[ 315] =  'sd12910;
    data[ 316] =  'sd64550;
    data[ 317] = -'sd4932;
    data[ 318] = -'sd24660;
    data[ 319] =  'sd40541;
    data[ 320] =  'sd38864;
    data[ 321] =  'sd30479;
    data[ 322] = -'sd11446;
    data[ 323] = -'sd57230;
    data[ 324] =  'sd41532;
    data[ 325] =  'sd43819;
    data[ 326] =  'sd55254;
    data[ 327] = -'sd51412;
    data[ 328] =  'sd70622;
    data[ 329] =  'sd25428;
    data[ 330] = -'sd36701;
    data[ 331] = -'sd19664;
    data[ 332] =  'sd65521;
    data[ 333] = -'sd77;
    data[ 334] = -'sd385;
    data[ 335] = -'sd1925;
    data[ 336] = -'sd9625;
    data[ 337] = -'sd48125;
    data[ 338] = -'sd76784;
    data[ 339] = -'sd56238;
    data[ 340] =  'sd46492;
    data[ 341] =  'sd68619;
    data[ 342] =  'sd15413;
    data[ 343] =  'sd77065;
    data[ 344] =  'sd57643;
    data[ 345] = -'sd39467;
    data[ 346] = -'sd33494;
    data[ 347] = -'sd3629;
    data[ 348] = -'sd18145;
    data[ 349] =  'sd73116;
    data[ 350] =  'sd37898;
    data[ 351] =  'sd25649;
    data[ 352] = -'sd35596;
    data[ 353] = -'sd14139;
    data[ 354] = -'sd70695;
    data[ 355] = -'sd25793;
    data[ 356] =  'sd34876;
    data[ 357] =  'sd10539;
    data[ 358] =  'sd52695;
    data[ 359] = -'sd64207;
    data[ 360] =  'sd6647;
    data[ 361] =  'sd33235;
    data[ 362] =  'sd2334;
    data[ 363] =  'sd11670;
    data[ 364] =  'sd58350;
    data[ 365] = -'sd35932;
    data[ 366] = -'sd15819;
    data[ 367] = -'sd79095;
    data[ 368] = -'sd67793;
    data[ 369] = -'sd11283;
    data[ 370] = -'sd56415;
    data[ 371] =  'sd45607;
    data[ 372] =  'sd64194;
    data[ 373] = -'sd6712;
    data[ 374] = -'sd33560;
    data[ 375] = -'sd3959;
    data[ 376] = -'sd19795;
    data[ 377] =  'sd64866;
    data[ 378] = -'sd3352;
    data[ 379] = -'sd16760;
    data[ 380] =  'sd80041;
    data[ 381] =  'sd72523;
    data[ 382] =  'sd34933;
    data[ 383] =  'sd10824;
    data[ 384] =  'sd54120;
    data[ 385] = -'sd57082;
    data[ 386] =  'sd42272;
    data[ 387] =  'sd47519;
    data[ 388] =  'sd73754;
    data[ 389] =  'sd41088;
    data[ 390] =  'sd41599;
    data[ 391] =  'sd44154;
    data[ 392] =  'sd56929;
    data[ 393] = -'sd43037;
    data[ 394] = -'sd51344;
    data[ 395] =  'sd70962;
    data[ 396] =  'sd27128;
    data[ 397] = -'sd28201;
    data[ 398] =  'sd22836;
    data[ 399] = -'sd49661;
    data[ 400] =  'sd79377;
    data[ 401] =  'sd69203;
    data[ 402] =  'sd18333;
    data[ 403] = -'sd72176;
    data[ 404] = -'sd33198;
    data[ 405] = -'sd2149;
    data[ 406] = -'sd10745;
    data[ 407] = -'sd53725;
    data[ 408] =  'sd59057;
    data[ 409] = -'sd32397;
    data[ 410] =  'sd1856;
    data[ 411] =  'sd9280;
    data[ 412] =  'sd46400;
    data[ 413] =  'sd68159;
    data[ 414] =  'sd13113;
    data[ 415] =  'sd65565;
    data[ 416] =  'sd143;
    data[ 417] =  'sd715;
    data[ 418] =  'sd3575;
    data[ 419] =  'sd17875;
    data[ 420] = -'sd74466;
    data[ 421] = -'sd44648;
    data[ 422] = -'sd59399;
    data[ 423] =  'sd30687;
    data[ 424] = -'sd10406;
    data[ 425] = -'sd52030;
    data[ 426] =  'sd67532;
    data[ 427] =  'sd9978;
    data[ 428] =  'sd49890;
    data[ 429] = -'sd78232;
    data[ 430] = -'sd63478;
    data[ 431] =  'sd10292;
    data[ 432] =  'sd51460;
    data[ 433] = -'sd70382;
    data[ 434] = -'sd24228;
    data[ 435] =  'sd42701;
    data[ 436] =  'sd49664;
    data[ 437] = -'sd79362;
    data[ 438] = -'sd69128;
    data[ 439] = -'sd17958;
    data[ 440] =  'sd74051;
    data[ 441] =  'sd42573;
    data[ 442] =  'sd49024;
    data[ 443] =  'sd81279;
    data[ 444] =  'sd78713;
    data[ 445] =  'sd65883;
    data[ 446] =  'sd1733;
    data[ 447] =  'sd8665;
    data[ 448] =  'sd43325;
    data[ 449] =  'sd52784;
    data[ 450] = -'sd63762;
    data[ 451] =  'sd8872;
    data[ 452] =  'sd44360;
    data[ 453] =  'sd57959;
    data[ 454] = -'sd37887;
    data[ 455] = -'sd25594;
    data[ 456] =  'sd35871;
    data[ 457] =  'sd15514;
    data[ 458] =  'sd77570;
    data[ 459] =  'sd60168;
    data[ 460] = -'sd26842;
    data[ 461] =  'sd29631;
    data[ 462] = -'sd15686;
    data[ 463] = -'sd78430;
    data[ 464] = -'sd64468;
    data[ 465] =  'sd5342;
    data[ 466] =  'sd26710;
    data[ 467] = -'sd30291;
    data[ 468] =  'sd12386;
    data[ 469] =  'sd61930;
    data[ 470] = -'sd18032;
    data[ 471] =  'sd73681;
    data[ 472] =  'sd40723;
    data[ 473] =  'sd39774;
    data[ 474] =  'sd35029;
    data[ 475] =  'sd11304;
    data[ 476] =  'sd56520;
    data[ 477] = -'sd45082;
    data[ 478] = -'sd61569;
    data[ 479] =  'sd19837;
    data[ 480] = -'sd64656;
    data[ 481] =  'sd4402;
    data[ 482] =  'sd22010;
    data[ 483] = -'sd53791;
    data[ 484] =  'sd58727;
    data[ 485] = -'sd34047;
    data[ 486] = -'sd6394;
    data[ 487] = -'sd31970;
    data[ 488] =  'sd3991;
    data[ 489] =  'sd19955;
    data[ 490] = -'sd64066;
    data[ 491] =  'sd7352;
    data[ 492] =  'sd36760;
    data[ 493] =  'sd19959;
    data[ 494] = -'sd64046;
    data[ 495] =  'sd7452;
    data[ 496] =  'sd37260;
    data[ 497] =  'sd22459;
    data[ 498] = -'sd51546;
    data[ 499] =  'sd69952;
    data[ 500] =  'sd22078;
    data[ 501] = -'sd53451;
    data[ 502] =  'sd60427;
    data[ 503] = -'sd25547;
    data[ 504] =  'sd36106;
    data[ 505] =  'sd16689;
    data[ 506] = -'sd80396;
    data[ 507] = -'sd74298;
    data[ 508] = -'sd43808;
    data[ 509] = -'sd55199;
    data[ 510] =  'sd51687;
    data[ 511] = -'sd69247;
    data[ 512] = -'sd18553;
    data[ 513] =  'sd71076;
    data[ 514] =  'sd27698;
    data[ 515] = -'sd25351;
    data[ 516] =  'sd37086;
    data[ 517] =  'sd21589;
    data[ 518] = -'sd55896;
    data[ 519] =  'sd48202;
    data[ 520] =  'sd77169;
    data[ 521] =  'sd58163;
    data[ 522] = -'sd36867;
    data[ 523] = -'sd20494;
    data[ 524] =  'sd61371;
    data[ 525] = -'sd20827;
    data[ 526] =  'sd59706;
    data[ 527] = -'sd29152;
    data[ 528] =  'sd18081;
    data[ 529] = -'sd73436;
    data[ 530] = -'sd39498;
    data[ 531] = -'sd33649;
    data[ 532] = -'sd4404;
    data[ 533] = -'sd22020;
    data[ 534] =  'sd53741;
    data[ 535] = -'sd58977;
    data[ 536] =  'sd32797;
    data[ 537] =  'sd144;
    data[ 538] =  'sd720;
    data[ 539] =  'sd3600;
    data[ 540] =  'sd18000;
    data[ 541] = -'sd73841;
    data[ 542] = -'sd41523;
    data[ 543] = -'sd43774;
    data[ 544] = -'sd55029;
    data[ 545] =  'sd52537;
    data[ 546] = -'sd64997;
    data[ 547] =  'sd2697;
    data[ 548] =  'sd13485;
    data[ 549] =  'sd67425;
    data[ 550] =  'sd9443;
    data[ 551] =  'sd47215;
    data[ 552] =  'sd72234;
    data[ 553] =  'sd33488;
    data[ 554] =  'sd3599;
    data[ 555] =  'sd17995;
    data[ 556] = -'sd73866;
    data[ 557] = -'sd41648;
    data[ 558] = -'sd44399;
    data[ 559] = -'sd58154;
    data[ 560] =  'sd36912;
    data[ 561] =  'sd20719;
    data[ 562] = -'sd60246;
    data[ 563] =  'sd26452;
    data[ 564] = -'sd31581;
    data[ 565] =  'sd5936;
    data[ 566] =  'sd29680;
    data[ 567] = -'sd15441;
    data[ 568] = -'sd77205;
    data[ 569] = -'sd58343;
    data[ 570] =  'sd35967;
    data[ 571] =  'sd15994;
    data[ 572] =  'sd79970;
    data[ 573] =  'sd72168;
    data[ 574] =  'sd33158;
    data[ 575] =  'sd1949;
    data[ 576] =  'sd9745;
    data[ 577] =  'sd48725;
    data[ 578] =  'sd79784;
    data[ 579] =  'sd71238;
    data[ 580] =  'sd28508;
    data[ 581] = -'sd21301;
    data[ 582] =  'sd57336;
    data[ 583] = -'sd41002;
    data[ 584] = -'sd41169;
    data[ 585] = -'sd42004;
    data[ 586] = -'sd46179;
    data[ 587] = -'sd67054;
    data[ 588] = -'sd7588;
    data[ 589] = -'sd37940;
    data[ 590] = -'sd25859;
    data[ 591] =  'sd34546;
    data[ 592] =  'sd8889;
    data[ 593] =  'sd44445;
    data[ 594] =  'sd58384;
    data[ 595] = -'sd35762;
    data[ 596] = -'sd14969;
    data[ 597] = -'sd74845;
    data[ 598] = -'sd46543;
    data[ 599] = -'sd68874;
    data[ 600] = -'sd16688;
    data[ 601] =  'sd80401;
    data[ 602] =  'sd74323;
    data[ 603] =  'sd43933;
    data[ 604] =  'sd55824;
    data[ 605] = -'sd48562;
    data[ 606] = -'sd78969;
    data[ 607] = -'sd67163;
    data[ 608] = -'sd8133;
    data[ 609] = -'sd40665;
    data[ 610] = -'sd39484;
    data[ 611] = -'sd33579;
    data[ 612] = -'sd4054;
    data[ 613] = -'sd20270;
    data[ 614] =  'sd62491;
    data[ 615] = -'sd15227;
    data[ 616] = -'sd76135;
    data[ 617] = -'sd52993;
    data[ 618] =  'sd62717;
    data[ 619] = -'sd14097;
    data[ 620] = -'sd70485;
    data[ 621] = -'sd24743;
    data[ 622] =  'sd40126;
    data[ 623] =  'sd36789;
    data[ 624] =  'sd20104;
    data[ 625] = -'sd63321;
    data[ 626] =  'sd11077;
    data[ 627] =  'sd55385;
    data[ 628] = -'sd50757;
    data[ 629] =  'sd73897;
    data[ 630] =  'sd41803;
    data[ 631] =  'sd45174;
    data[ 632] =  'sd62029;
    data[ 633] = -'sd17537;
    data[ 634] =  'sd76156;
    data[ 635] =  'sd53098;
    data[ 636] = -'sd62192;
    data[ 637] =  'sd16722;
    data[ 638] = -'sd80231;
    data[ 639] = -'sd73473;
    data[ 640] = -'sd39683;
    data[ 641] = -'sd34574;
    data[ 642] = -'sd9029;
    data[ 643] = -'sd45145;
    data[ 644] = -'sd61884;
    data[ 645] =  'sd18262;
    data[ 646] = -'sd72531;
    data[ 647] = -'sd34973;
    data[ 648] = -'sd11024;
    data[ 649] = -'sd55120;
    data[ 650] =  'sd52082;
    data[ 651] = -'sd67272;
    data[ 652] = -'sd8678;
    data[ 653] = -'sd43390;
    data[ 654] = -'sd53109;
    data[ 655] =  'sd62137;
    data[ 656] = -'sd16997;
    data[ 657] =  'sd78856;
    data[ 658] =  'sd66598;
    data[ 659] =  'sd5308;
    data[ 660] =  'sd26540;
    data[ 661] = -'sd31141;
    data[ 662] =  'sd8136;
    data[ 663] =  'sd40680;
    data[ 664] =  'sd39559;
    data[ 665] =  'sd33954;
    data[ 666] =  'sd5929;
    data[ 667] =  'sd29645;
    data[ 668] = -'sd15616;
    data[ 669] = -'sd78080;
    data[ 670] = -'sd62718;
    data[ 671] =  'sd14092;
    data[ 672] =  'sd70460;
    data[ 673] =  'sd24618;
    data[ 674] = -'sd40751;
    data[ 675] = -'sd39914;
    data[ 676] = -'sd35729;
    data[ 677] = -'sd14804;
    data[ 678] = -'sd74020;
    data[ 679] = -'sd42418;
    data[ 680] = -'sd48249;
    data[ 681] = -'sd77404;
    data[ 682] = -'sd59338;
    data[ 683] =  'sd30992;
    data[ 684] = -'sd8881;
    data[ 685] = -'sd44405;
    data[ 686] = -'sd58184;
    data[ 687] =  'sd36762;
    data[ 688] =  'sd19969;
    data[ 689] = -'sd63996;
    data[ 690] =  'sd7702;
    data[ 691] =  'sd38510;
    data[ 692] =  'sd28709;
    data[ 693] = -'sd20296;
    data[ 694] =  'sd62361;
    data[ 695] = -'sd15877;
    data[ 696] = -'sd79385;
    data[ 697] = -'sd69243;
    data[ 698] = -'sd18533;
    data[ 699] =  'sd71176;
    data[ 700] =  'sd28198;
    data[ 701] = -'sd22851;
    data[ 702] =  'sd49586;
    data[ 703] = -'sd79752;
    data[ 704] = -'sd71078;
    data[ 705] = -'sd27708;
    data[ 706] =  'sd25301;
    data[ 707] = -'sd37336;
    data[ 708] = -'sd22839;
    data[ 709] =  'sd49646;
    data[ 710] = -'sd79452;
    data[ 711] = -'sd69578;
    data[ 712] = -'sd20208;
    data[ 713] =  'sd62801;
    data[ 714] = -'sd13677;
    data[ 715] = -'sd68385;
    data[ 716] = -'sd14243;
    data[ 717] = -'sd71215;
    data[ 718] = -'sd28393;
    data[ 719] =  'sd21876;
    data[ 720] = -'sd54461;
    data[ 721] =  'sd55377;
    data[ 722] = -'sd50797;
    data[ 723] =  'sd73697;
    data[ 724] =  'sd40803;
    data[ 725] =  'sd40174;
    data[ 726] =  'sd37029;
    data[ 727] =  'sd21304;
    data[ 728] = -'sd57321;
    data[ 729] =  'sd41077;
    data[ 730] =  'sd41544;
    data[ 731] =  'sd43879;
    data[ 732] =  'sd55554;
    data[ 733] = -'sd49912;
    data[ 734] =  'sd78122;
    data[ 735] =  'sd62928;
    data[ 736] = -'sd13042;
    data[ 737] = -'sd65210;
    data[ 738] =  'sd1632;
    data[ 739] =  'sd8160;
    data[ 740] =  'sd40800;
    data[ 741] =  'sd40159;
    data[ 742] =  'sd36954;
    data[ 743] =  'sd20929;
    data[ 744] = -'sd59196;
    data[ 745] =  'sd31702;
    data[ 746] = -'sd5331;
    data[ 747] = -'sd26655;
    data[ 748] =  'sd30566;
    data[ 749] = -'sd11011;
    data[ 750] = -'sd55055;
    data[ 751] =  'sd52407;
    data[ 752] = -'sd65647;
    data[ 753] = -'sd553;
    data[ 754] = -'sd2765;
    data[ 755] = -'sd13825;
    data[ 756] = -'sd69125;
    data[ 757] = -'sd17943;
    data[ 758] =  'sd74126;
    data[ 759] =  'sd42948;
    data[ 760] =  'sd50899;
    data[ 761] = -'sd73187;
    data[ 762] = -'sd38253;
    data[ 763] = -'sd27424;
    data[ 764] =  'sd26721;
    data[ 765] = -'sd30236;
    data[ 766] =  'sd12661;
    data[ 767] =  'sd63305;
    data[ 768] = -'sd11157;
    data[ 769] = -'sd55785;
    data[ 770] =  'sd48757;
    data[ 771] =  'sd79944;
    data[ 772] =  'sd72038;
    data[ 773] =  'sd32508;
    data[ 774] = -'sd1301;
    data[ 775] = -'sd6505;
    data[ 776] = -'sd32525;
    data[ 777] =  'sd1216;
    data[ 778] =  'sd6080;
    data[ 779] =  'sd30400;
    data[ 780] = -'sd11841;
    data[ 781] = -'sd59205;
    data[ 782] =  'sd31657;
    data[ 783] = -'sd5556;
    data[ 784] = -'sd27780;
    data[ 785] =  'sd24941;
    data[ 786] = -'sd39136;
    data[ 787] = -'sd31839;
    data[ 788] =  'sd4646;
    data[ 789] =  'sd23230;
    data[ 790] = -'sd47691;
    data[ 791] = -'sd74614;
    data[ 792] = -'sd45388;
    data[ 793] = -'sd63099;
    data[ 794] =  'sd12187;
    data[ 795] =  'sd60935;
    data[ 796] = -'sd23007;
    data[ 797] =  'sd48806;
    data[ 798] =  'sd80189;
    data[ 799] =  'sd73263;
    data[ 800] =  'sd38633;
    data[ 801] =  'sd29324;
    data[ 802] = -'sd17221;
    data[ 803] =  'sd77736;
    data[ 804] =  'sd60998;
    data[ 805] = -'sd22692;
    data[ 806] =  'sd50381;
    data[ 807] = -'sd75777;
    data[ 808] = -'sd51203;
    data[ 809] =  'sd71667;
    data[ 810] =  'sd30653;
    data[ 811] = -'sd10576;
    data[ 812] = -'sd52880;
    data[ 813] =  'sd63282;
    data[ 814] = -'sd11272;
    data[ 815] = -'sd56360;
    data[ 816] =  'sd45882;
    data[ 817] =  'sd65569;
    data[ 818] =  'sd163;
    data[ 819] =  'sd815;
    data[ 820] =  'sd4075;
    data[ 821] =  'sd20375;
    data[ 822] = -'sd61966;
    data[ 823] =  'sd17852;
    data[ 824] = -'sd74581;
    data[ 825] = -'sd45223;
    data[ 826] = -'sd62274;
    data[ 827] =  'sd16312;
    data[ 828] =  'sd81560;
    data[ 829] =  'sd80118;
    data[ 830] =  'sd72908;
    data[ 831] =  'sd36858;
    data[ 832] =  'sd20449;
    data[ 833] = -'sd61596;
    data[ 834] =  'sd19702;
    data[ 835] = -'sd65331;
    data[ 836] =  'sd1027;
    data[ 837] =  'sd5135;
    data[ 838] =  'sd25675;
    data[ 839] = -'sd35466;
    data[ 840] = -'sd13489;
    data[ 841] = -'sd67445;
    data[ 842] = -'sd9543;
    data[ 843] = -'sd47715;
    data[ 844] = -'sd74734;
    data[ 845] = -'sd45988;
    data[ 846] = -'sd66099;
    data[ 847] = -'sd2813;
    data[ 848] = -'sd14065;
    data[ 849] = -'sd70325;
    data[ 850] = -'sd23943;
    data[ 851] =  'sd44126;
    data[ 852] =  'sd56789;
    data[ 853] = -'sd43737;
    data[ 854] = -'sd54844;
    data[ 855] =  'sd53462;
    data[ 856] = -'sd60372;
    data[ 857] =  'sd25822;
    data[ 858] = -'sd34731;
    data[ 859] = -'sd9814;
    data[ 860] = -'sd49070;
    data[ 861] = -'sd81509;
    data[ 862] = -'sd79863;
    data[ 863] = -'sd71633;
    data[ 864] = -'sd30483;
    data[ 865] =  'sd11426;
    data[ 866] =  'sd57130;
    data[ 867] = -'sd42032;
    data[ 868] = -'sd46319;
    data[ 869] = -'sd67754;
    data[ 870] = -'sd11088;
    data[ 871] = -'sd55440;
    data[ 872] =  'sd50482;
    data[ 873] = -'sd75272;
    data[ 874] = -'sd48678;
    data[ 875] = -'sd79549;
    data[ 876] = -'sd70063;
    data[ 877] = -'sd22633;
    data[ 878] =  'sd50676;
    data[ 879] = -'sd74302;
    data[ 880] = -'sd43828;
    data[ 881] = -'sd55299;
    data[ 882] =  'sd51187;
    data[ 883] = -'sd71747;
    data[ 884] = -'sd31053;
    data[ 885] =  'sd8576;
    data[ 886] =  'sd42880;
    data[ 887] =  'sd50559;
    data[ 888] = -'sd74887;
    data[ 889] = -'sd46753;
    data[ 890] = -'sd69924;
    data[ 891] = -'sd21938;
    data[ 892] =  'sd54151;
    data[ 893] = -'sd56927;
    data[ 894] =  'sd43047;
    data[ 895] =  'sd51394;
    data[ 896] = -'sd70712;
    data[ 897] = -'sd25878;
    data[ 898] =  'sd34451;
    data[ 899] =  'sd8414;
    data[ 900] =  'sd42070;
    data[ 901] =  'sd46509;
    data[ 902] =  'sd68704;
    data[ 903] =  'sd15838;
    data[ 904] =  'sd79190;
    data[ 905] =  'sd68268;
    data[ 906] =  'sd13658;
    data[ 907] =  'sd68290;
    data[ 908] =  'sd13768;
    data[ 909] =  'sd68840;
    data[ 910] =  'sd16518;
    data[ 911] = -'sd81251;
    data[ 912] = -'sd78573;
    data[ 913] = -'sd65183;
    data[ 914] =  'sd1767;
    data[ 915] =  'sd8835;
    data[ 916] =  'sd44175;
    data[ 917] =  'sd57034;
    data[ 918] = -'sd42512;
    data[ 919] = -'sd48719;
    data[ 920] = -'sd79754;
    data[ 921] = -'sd71088;
    data[ 922] = -'sd27758;
    data[ 923] =  'sd25051;
    data[ 924] = -'sd38586;
    data[ 925] = -'sd29089;
    data[ 926] =  'sd18396;
    data[ 927] = -'sd71861;
    data[ 928] = -'sd31623;
    data[ 929] =  'sd5726;
    data[ 930] =  'sd28630;
    data[ 931] = -'sd20691;
    data[ 932] =  'sd60386;
    data[ 933] = -'sd25752;
    data[ 934] =  'sd35081;
    data[ 935] =  'sd11564;
    data[ 936] =  'sd57820;
    data[ 937] = -'sd38582;
    data[ 938] = -'sd29069;
    data[ 939] =  'sd18496;
    data[ 940] = -'sd71361;
    data[ 941] = -'sd29123;
    data[ 942] =  'sd18226;
    data[ 943] = -'sd72711;
    data[ 944] = -'sd35873;
    data[ 945] = -'sd15524;
    data[ 946] = -'sd77620;
    data[ 947] = -'sd60418;
    data[ 948] =  'sd25592;
    data[ 949] = -'sd35881;
    data[ 950] = -'sd15564;
    data[ 951] = -'sd77820;
    data[ 952] = -'sd61418;
    data[ 953] =  'sd20592;
    data[ 954] = -'sd60881;
    data[ 955] =  'sd23277;
    data[ 956] = -'sd47456;
    data[ 957] = -'sd73439;
    data[ 958] = -'sd39513;
    data[ 959] = -'sd33724;
    data[ 960] = -'sd4779;
    data[ 961] = -'sd23895;
    data[ 962] =  'sd44366;
    data[ 963] =  'sd57989;
    data[ 964] = -'sd37737;
    data[ 965] = -'sd24844;
    data[ 966] =  'sd39621;
    data[ 967] =  'sd34264;
    data[ 968] =  'sd7479;
    data[ 969] =  'sd37395;
    data[ 970] =  'sd23134;
    data[ 971] = -'sd48171;
    data[ 972] = -'sd77014;
    data[ 973] = -'sd57388;
    data[ 974] =  'sd40742;
    data[ 975] =  'sd39869;
    data[ 976] =  'sd35504;
    data[ 977] =  'sd13679;
    data[ 978] =  'sd68395;
    data[ 979] =  'sd14293;
    data[ 980] =  'sd71465;
    data[ 981] =  'sd29643;
    data[ 982] = -'sd15626;
    data[ 983] = -'sd78130;
    data[ 984] = -'sd62968;
    data[ 985] =  'sd12842;
    data[ 986] =  'sd64210;
    data[ 987] = -'sd6632;
    data[ 988] = -'sd33160;
    data[ 989] = -'sd1959;
    data[ 990] = -'sd9795;
    data[ 991] = -'sd48975;
    data[ 992] = -'sd81034;
    data[ 993] = -'sd77488;
    data[ 994] = -'sd59758;
    data[ 995] =  'sd28892;
    data[ 996] = -'sd19381;
    data[ 997] =  'sd66936;
    data[ 998] =  'sd6998;
    data[ 999] =  'sd34990;
    data[1000] =  'sd11109;
    data[1001] =  'sd55545;
    data[1002] = -'sd49957;
    data[1003] =  'sd77897;
    data[1004] =  'sd61803;
    data[1005] = -'sd18667;
    data[1006] =  'sd70506;
    data[1007] =  'sd24848;
    data[1008] = -'sd39601;
    data[1009] = -'sd34164;
    data[1010] = -'sd6979;
    data[1011] = -'sd34895;
    data[1012] = -'sd10634;
    data[1013] = -'sd53170;
    data[1014] =  'sd61832;
    data[1015] = -'sd18522;
    data[1016] =  'sd71231;
    data[1017] =  'sd28473;
    data[1018] = -'sd21476;
    data[1019] =  'sd56461;
    data[1020] = -'sd45377;
    data[1021] = -'sd63044;
    data[1022] =  'sd12462;
    data[1023] =  'sd62310;
    data[1024] = -'sd16132;
    data[1025] = -'sd80660;
    data[1026] = -'sd75618;
    data[1027] = -'sd50408;
    data[1028] =  'sd75642;
    data[1029] =  'sd50528;
    data[1030] = -'sd75042;
    data[1031] = -'sd47528;
    data[1032] = -'sd73799;
    data[1033] = -'sd41313;
    data[1034] = -'sd42724;
    data[1035] = -'sd49779;
    data[1036] =  'sd78787;
    data[1037] =  'sd66253;
    data[1038] =  'sd3583;
    data[1039] =  'sd17915;
    data[1040] = -'sd74266;
    data[1041] = -'sd43648;
    data[1042] = -'sd54399;
    data[1043] =  'sd55687;
    data[1044] = -'sd49247;
    data[1045] =  'sd81447;
    data[1046] =  'sd79553;
    data[1047] =  'sd70083;
    data[1048] =  'sd22733;
    data[1049] = -'sd50176;
    data[1050] =  'sd76802;
    data[1051] =  'sd56328;
    data[1052] = -'sd46042;
    data[1053] = -'sd66369;
    data[1054] = -'sd4163;
    data[1055] = -'sd20815;
    data[1056] =  'sd59766;
    data[1057] = -'sd28852;
    data[1058] =  'sd19581;
    data[1059] = -'sd65936;
    data[1060] = -'sd1998;
    data[1061] = -'sd9990;
    data[1062] = -'sd49950;
    data[1063] =  'sd77932;
    data[1064] =  'sd61978;
    data[1065] = -'sd17792;
    data[1066] =  'sd74881;
    data[1067] =  'sd46723;
    data[1068] =  'sd69774;
    data[1069] =  'sd21188;
    data[1070] = -'sd57901;
    data[1071] =  'sd38177;
    data[1072] =  'sd27044;
    data[1073] = -'sd28621;
    data[1074] =  'sd20736;
    data[1075] = -'sd60161;
    data[1076] =  'sd26877;
    data[1077] = -'sd29456;
    data[1078] =  'sd16561;
    data[1079] = -'sd81036;
    data[1080] = -'sd77498;
    data[1081] = -'sd59808;
    data[1082] =  'sd28642;
    data[1083] = -'sd20631;
    data[1084] =  'sd60686;
    data[1085] = -'sd24252;
    data[1086] =  'sd42581;
    data[1087] =  'sd49064;
    data[1088] =  'sd81479;
    data[1089] =  'sd79713;
    data[1090] =  'sd70883;
    data[1091] =  'sd26733;
    data[1092] = -'sd30176;
    data[1093] =  'sd12961;
    data[1094] =  'sd64805;
    data[1095] = -'sd3657;
    data[1096] = -'sd18285;
    data[1097] =  'sd72416;
    data[1098] =  'sd34398;
    data[1099] =  'sd8149;
    data[1100] =  'sd40745;
    data[1101] =  'sd39884;
    data[1102] =  'sd35579;
    data[1103] =  'sd14054;
    data[1104] =  'sd70270;
    data[1105] =  'sd23668;
    data[1106] = -'sd45501;
    data[1107] = -'sd63664;
    data[1108] =  'sd9362;
    data[1109] =  'sd46810;
    data[1110] =  'sd70209;
    data[1111] =  'sd23363;
    data[1112] = -'sd47026;
    data[1113] = -'sd71289;
    data[1114] = -'sd28763;
    data[1115] =  'sd20026;
    data[1116] = -'sd63711;
    data[1117] =  'sd9127;
    data[1118] =  'sd45635;
    data[1119] =  'sd64334;
    data[1120] = -'sd6012;
    data[1121] = -'sd30060;
    data[1122] =  'sd13541;
    data[1123] =  'sd67705;
    data[1124] =  'sd10843;
    data[1125] =  'sd54215;
    data[1126] = -'sd56607;
    data[1127] =  'sd44647;
    data[1128] =  'sd59394;
    data[1129] = -'sd30712;
    data[1130] =  'sd10281;
    data[1131] =  'sd51405;
    data[1132] = -'sd70657;
    data[1133] = -'sd25603;
    data[1134] =  'sd35826;
    data[1135] =  'sd15289;
    data[1136] =  'sd76445;
    data[1137] =  'sd54543;
    data[1138] = -'sd54967;
    data[1139] =  'sd52847;
    data[1140] = -'sd63447;
    data[1141] =  'sd10447;
    data[1142] =  'sd52235;
    data[1143] = -'sd66507;
    data[1144] = -'sd4853;
    data[1145] = -'sd24265;
    data[1146] =  'sd42516;
    data[1147] =  'sd48739;
    data[1148] =  'sd79854;
    data[1149] =  'sd71588;
    data[1150] =  'sd30258;
    data[1151] = -'sd12551;
    data[1152] = -'sd62755;
    data[1153] =  'sd13907;
    data[1154] =  'sd69535;
    data[1155] =  'sd19993;
    data[1156] = -'sd63876;
    data[1157] =  'sd8302;
    data[1158] =  'sd41510;
    data[1159] =  'sd43709;
    data[1160] =  'sd54704;
    data[1161] = -'sd54162;
    data[1162] =  'sd56872;
    data[1163] = -'sd43322;
    data[1164] = -'sd52769;
    data[1165] =  'sd63837;
    data[1166] = -'sd8497;
    data[1167] = -'sd42485;
    data[1168] = -'sd48584;
    data[1169] = -'sd79079;
    data[1170] = -'sd67713;
    data[1171] = -'sd10883;
    data[1172] = -'sd54415;
    data[1173] =  'sd55607;
    data[1174] = -'sd49647;
    data[1175] =  'sd79447;
    data[1176] =  'sd69553;
    data[1177] =  'sd20083;
    data[1178] = -'sd63426;
    data[1179] =  'sd10552;
    data[1180] =  'sd52760;
    data[1181] = -'sd63882;
    data[1182] =  'sd8272;
    data[1183] =  'sd41360;
    data[1184] =  'sd42959;
    data[1185] =  'sd50954;
    data[1186] = -'sd72912;
    data[1187] = -'sd36878;
    data[1188] = -'sd20549;
    data[1189] =  'sd61096;
    data[1190] = -'sd22202;
    data[1191] =  'sd52831;
    data[1192] = -'sd63527;
    data[1193] =  'sd10047;
    data[1194] =  'sd50235;
    data[1195] = -'sd76507;
    data[1196] = -'sd54853;
    data[1197] =  'sd53417;
    data[1198] = -'sd60597;
    data[1199] =  'sd24697;
    data[1200] = -'sd40356;
    data[1201] = -'sd37939;
    data[1202] = -'sd25854;
    data[1203] =  'sd34571;
    data[1204] =  'sd9014;
    data[1205] =  'sd45070;
    data[1206] =  'sd61509;
    data[1207] = -'sd20137;
    data[1208] =  'sd63156;
    data[1209] = -'sd11902;
    data[1210] = -'sd59510;
    data[1211] =  'sd30132;
    data[1212] = -'sd13181;
    data[1213] = -'sd65905;
    data[1214] = -'sd1843;
    data[1215] = -'sd9215;
    data[1216] = -'sd46075;
    data[1217] = -'sd66534;
    data[1218] = -'sd4988;
    data[1219] = -'sd24940;
    data[1220] =  'sd39141;
    data[1221] =  'sd31864;
    data[1222] = -'sd4521;
    data[1223] = -'sd22605;
    data[1224] =  'sd50816;
    data[1225] = -'sd73602;
    data[1226] = -'sd40328;
    data[1227] = -'sd37799;
    data[1228] = -'sd25154;
    data[1229] =  'sd38071;
    data[1230] =  'sd26514;
    data[1231] = -'sd31271;
    data[1232] =  'sd7486;
    data[1233] =  'sd37430;
    data[1234] =  'sd23309;
    data[1235] = -'sd47296;
    data[1236] = -'sd72639;
    data[1237] = -'sd35513;
    data[1238] = -'sd13724;
    data[1239] = -'sd68620;
    data[1240] = -'sd15418;
    data[1241] = -'sd77090;
    data[1242] = -'sd57768;
    data[1243] =  'sd38842;
    data[1244] =  'sd30369;
    data[1245] = -'sd11996;
    data[1246] = -'sd59980;
    data[1247] =  'sd27782;
    data[1248] = -'sd24931;
    data[1249] =  'sd39186;
    data[1250] =  'sd32089;
    data[1251] = -'sd3396;
    data[1252] = -'sd16980;
    data[1253] =  'sd78941;
    data[1254] =  'sd67023;
    data[1255] =  'sd7433;
    data[1256] =  'sd37165;
    data[1257] =  'sd21984;
    data[1258] = -'sd53921;
    data[1259] =  'sd58077;
    data[1260] = -'sd37297;
    data[1261] = -'sd22644;
    data[1262] =  'sd50621;
    data[1263] = -'sd74577;
    data[1264] = -'sd45203;
    data[1265] = -'sd62174;
    data[1266] =  'sd16812;
    data[1267] = -'sd79781;
    data[1268] = -'sd71223;
    data[1269] = -'sd28433;
    data[1270] =  'sd21676;
    data[1271] = -'sd55461;
    data[1272] =  'sd50377;
    data[1273] = -'sd75797;
    data[1274] = -'sd51303;
    data[1275] =  'sd71167;
    data[1276] =  'sd28153;
    data[1277] = -'sd23076;
    data[1278] =  'sd48461;
    data[1279] =  'sd78464;
    data[1280] =  'sd64638;
    data[1281] = -'sd4492;
    data[1282] = -'sd22460;
    data[1283] =  'sd51541;
    data[1284] = -'sd69977;
    data[1285] = -'sd22203;
    data[1286] =  'sd52826;
    data[1287] = -'sd63552;
    data[1288] =  'sd9922;
    data[1289] =  'sd49610;
    data[1290] = -'sd79632;
    data[1291] = -'sd70478;
    data[1292] = -'sd24708;
    data[1293] =  'sd40301;
    data[1294] =  'sd37664;
    data[1295] =  'sd24479;
    data[1296] = -'sd41446;
    data[1297] = -'sd43389;
    data[1298] = -'sd53104;
    data[1299] =  'sd62162;
    data[1300] = -'sd16872;
    data[1301] =  'sd79481;
    data[1302] =  'sd69723;
    data[1303] =  'sd20933;
    data[1304] = -'sd59176;
    data[1305] =  'sd31802;
    data[1306] = -'sd4831;
    data[1307] = -'sd24155;
    data[1308] =  'sd43066;
    data[1309] =  'sd51489;
    data[1310] = -'sd70237;
    data[1311] = -'sd23503;
    data[1312] =  'sd46326;
    data[1313] =  'sd67789;
    data[1314] =  'sd11263;
    data[1315] =  'sd56315;
    data[1316] = -'sd46107;
    data[1317] = -'sd66694;
    data[1318] = -'sd5788;
    data[1319] = -'sd28940;
    data[1320] =  'sd19141;
    data[1321] = -'sd68136;
    data[1322] = -'sd12998;
    data[1323] = -'sd64990;
    data[1324] =  'sd2732;
    data[1325] =  'sd13660;
    data[1326] =  'sd68300;
    data[1327] =  'sd13818;
    data[1328] =  'sd69090;
    data[1329] =  'sd17768;
    data[1330] = -'sd75001;
    data[1331] = -'sd47323;
    data[1332] = -'sd72774;
    data[1333] = -'sd36188;
    data[1334] = -'sd17099;
    data[1335] =  'sd78346;
    data[1336] =  'sd64048;
    data[1337] = -'sd7442;
    data[1338] = -'sd37210;
    data[1339] = -'sd22209;
    data[1340] =  'sd52796;
    data[1341] = -'sd63702;
    data[1342] =  'sd9172;
    data[1343] =  'sd45860;
    data[1344] =  'sd65459;
    data[1345] = -'sd387;
    data[1346] = -'sd1935;
    data[1347] = -'sd9675;
    data[1348] = -'sd48375;
    data[1349] = -'sd78034;
    data[1350] = -'sd62488;
    data[1351] =  'sd15242;
    data[1352] =  'sd76210;
    data[1353] =  'sd53368;
    data[1354] = -'sd60842;
    data[1355] =  'sd23472;
    data[1356] = -'sd46481;
    data[1357] = -'sd68564;
    data[1358] = -'sd15138;
    data[1359] = -'sd75690;
    data[1360] = -'sd50768;
    data[1361] =  'sd73842;
    data[1362] =  'sd41528;
    data[1363] =  'sd43799;
    data[1364] =  'sd55154;
    data[1365] = -'sd51912;
    data[1366] =  'sd68122;
    data[1367] =  'sd12928;
    data[1368] =  'sd64640;
    data[1369] = -'sd4482;
    data[1370] = -'sd22410;
    data[1371] =  'sd51791;
    data[1372] = -'sd68727;
    data[1373] = -'sd15953;
    data[1374] = -'sd79765;
    data[1375] = -'sd71143;
    data[1376] = -'sd28033;
    data[1377] =  'sd23676;
    data[1378] = -'sd45461;
    data[1379] = -'sd63464;
    data[1380] =  'sd10362;
    data[1381] =  'sd51810;
    data[1382] = -'sd68632;
    data[1383] = -'sd15478;
    data[1384] = -'sd77390;
    data[1385] = -'sd59268;
    data[1386] =  'sd31342;
    data[1387] = -'sd7131;
    data[1388] = -'sd35655;
    data[1389] = -'sd14434;
    data[1390] = -'sd72170;
    data[1391] = -'sd33168;
    data[1392] = -'sd1999;
    data[1393] = -'sd9995;
    data[1394] = -'sd49975;
    data[1395] =  'sd77807;
    data[1396] =  'sd61353;
    data[1397] = -'sd20917;
    data[1398] =  'sd59256;
    data[1399] = -'sd31402;
    data[1400] =  'sd6831;
    data[1401] =  'sd34155;
    data[1402] =  'sd6934;
    data[1403] =  'sd34670;
    data[1404] =  'sd9509;
    data[1405] =  'sd47545;
    data[1406] =  'sd73884;
    data[1407] =  'sd41738;
    data[1408] =  'sd44849;
    data[1409] =  'sd60404;
    data[1410] = -'sd25662;
    data[1411] =  'sd35531;
    data[1412] =  'sd13814;
    data[1413] =  'sd69070;
    data[1414] =  'sd17668;
    data[1415] = -'sd75501;
    data[1416] = -'sd49823;
    data[1417] =  'sd78567;
    data[1418] =  'sd65153;
    data[1419] = -'sd1917;
    data[1420] = -'sd9585;
    data[1421] = -'sd47925;
    data[1422] = -'sd75784;
    data[1423] = -'sd51238;
    data[1424] =  'sd71492;
    data[1425] =  'sd29778;
    data[1426] = -'sd14951;
    data[1427] = -'sd74755;
    data[1428] = -'sd46093;
    data[1429] = -'sd66624;
    data[1430] = -'sd5438;
    data[1431] = -'sd27190;
    data[1432] =  'sd27891;
    data[1433] = -'sd24386;
    data[1434] =  'sd41911;
    data[1435] =  'sd45714;
    data[1436] =  'sd64729;
    data[1437] = -'sd4037;
    data[1438] = -'sd20185;
    data[1439] =  'sd62916;
    data[1440] = -'sd13102;
    data[1441] = -'sd65510;
    data[1442] =  'sd132;
    data[1443] =  'sd660;
    data[1444] =  'sd3300;
    data[1445] =  'sd16500;
    data[1446] = -'sd81341;
    data[1447] = -'sd79023;
    data[1448] = -'sd67433;
    data[1449] = -'sd9483;
    data[1450] = -'sd47415;
    data[1451] = -'sd73234;
    data[1452] = -'sd38488;
    data[1453] = -'sd28599;
    data[1454] =  'sd20846;
    data[1455] = -'sd59611;
    data[1456] =  'sd29627;
    data[1457] = -'sd15706;
    data[1458] = -'sd78530;
    data[1459] = -'sd64968;
    data[1460] =  'sd2842;
    data[1461] =  'sd14210;
    data[1462] =  'sd71050;
    data[1463] =  'sd27568;
    data[1464] = -'sd26001;
    data[1465] =  'sd33836;
    data[1466] =  'sd5339;
    data[1467] =  'sd26695;
    data[1468] = -'sd30366;
    data[1469] =  'sd12011;
    data[1470] =  'sd60055;
    data[1471] = -'sd27407;
    data[1472] =  'sd26806;
    data[1473] = -'sd29811;
    data[1474] =  'sd14786;
    data[1475] =  'sd73930;
    data[1476] =  'sd41968;
    data[1477] =  'sd45999;
    data[1478] =  'sd66154;
    data[1479] =  'sd3088;
    data[1480] =  'sd15440;
    data[1481] =  'sd77200;
    data[1482] =  'sd58318;
    data[1483] = -'sd36092;
    data[1484] = -'sd16619;
    data[1485] =  'sd80746;
    data[1486] =  'sd76048;
    data[1487] =  'sd52558;
    data[1488] = -'sd64892;
    data[1489] =  'sd3222;
    data[1490] =  'sd16110;
    data[1491] =  'sd80550;
    data[1492] =  'sd75068;
    data[1493] =  'sd47658;
    data[1494] =  'sd74449;
    data[1495] =  'sd44563;
    data[1496] =  'sd58974;
    data[1497] = -'sd32812;
    data[1498] = -'sd219;
    data[1499] = -'sd1095;
    data[1500] = -'sd5475;
    data[1501] = -'sd27375;
    data[1502] =  'sd26966;
    data[1503] = -'sd29011;
    data[1504] =  'sd18786;
    data[1505] = -'sd69911;
    data[1506] = -'sd21873;
    data[1507] =  'sd54476;
    data[1508] = -'sd55302;
    data[1509] =  'sd51172;
    data[1510] = -'sd71822;
    data[1511] = -'sd31428;
    data[1512] =  'sd6701;
    data[1513] =  'sd33505;
    data[1514] =  'sd3684;
    data[1515] =  'sd18420;
    data[1516] = -'sd71741;
    data[1517] = -'sd31023;
    data[1518] =  'sd8726;
    data[1519] =  'sd43630;
    data[1520] =  'sd54309;
    data[1521] = -'sd56137;
    data[1522] =  'sd46997;
    data[1523] =  'sd71144;
    data[1524] =  'sd28038;
    data[1525] = -'sd23651;
    data[1526] =  'sd45586;
    data[1527] =  'sd64089;
    data[1528] = -'sd7237;
    data[1529] = -'sd36185;
    data[1530] = -'sd17084;
    data[1531] =  'sd78421;
    data[1532] =  'sd64423;
    data[1533] = -'sd5567;
    data[1534] = -'sd27835;
    data[1535] =  'sd24666;
    data[1536] = -'sd40511;
    data[1537] = -'sd38714;
    data[1538] = -'sd29729;
    data[1539] =  'sd15196;
    data[1540] =  'sd75980;
    data[1541] =  'sd52218;
    data[1542] = -'sd66592;
    data[1543] = -'sd5278;
    data[1544] = -'sd26390;
    data[1545] =  'sd31891;
    data[1546] = -'sd4386;
    data[1547] = -'sd21930;
    data[1548] =  'sd54191;
    data[1549] = -'sd56727;
    data[1550] =  'sd44047;
    data[1551] =  'sd56394;
    data[1552] = -'sd45712;
    data[1553] = -'sd64719;
    data[1554] =  'sd4087;
    data[1555] =  'sd20435;
    data[1556] = -'sd61666;
    data[1557] =  'sd19352;
    data[1558] = -'sd67081;
    data[1559] = -'sd7723;
    data[1560] = -'sd38615;
    data[1561] = -'sd29234;
    data[1562] =  'sd17671;
    data[1563] = -'sd75486;
    data[1564] = -'sd49748;
    data[1565] =  'sd78942;
    data[1566] =  'sd67028;
    data[1567] =  'sd7458;
    data[1568] =  'sd37290;
    data[1569] =  'sd22609;
    data[1570] = -'sd50796;
    data[1571] =  'sd73702;
    data[1572] =  'sd40828;
    data[1573] =  'sd40299;
    data[1574] =  'sd37654;
    data[1575] =  'sd24429;
    data[1576] = -'sd41696;
    data[1577] = -'sd44639;
    data[1578] = -'sd59354;
    data[1579] =  'sd30912;
    data[1580] = -'sd9281;
    data[1581] = -'sd46405;
    data[1582] = -'sd68184;
    data[1583] = -'sd13238;
    data[1584] = -'sd66190;
    data[1585] = -'sd3268;
    data[1586] = -'sd16340;
    data[1587] = -'sd81700;
    data[1588] = -'sd80818;
    data[1589] = -'sd76408;
    data[1590] = -'sd54358;
    data[1591] =  'sd55892;
    data[1592] = -'sd48222;
    data[1593] = -'sd77269;
    data[1594] = -'sd58663;
    data[1595] =  'sd34367;
    data[1596] =  'sd7994;
    data[1597] =  'sd39970;
    data[1598] =  'sd36009;
    data[1599] =  'sd16204;
    data[1600] =  'sd81020;
    data[1601] =  'sd77418;
    data[1602] =  'sd59408;
    data[1603] = -'sd30642;
    data[1604] =  'sd10631;
    data[1605] =  'sd53155;
    data[1606] = -'sd61907;
    data[1607] =  'sd18147;
    data[1608] = -'sd73106;
    data[1609] = -'sd37848;
    data[1610] = -'sd25399;
    data[1611] =  'sd36846;
    data[1612] =  'sd20389;
    data[1613] = -'sd61896;
    data[1614] =  'sd18202;
    data[1615] = -'sd72831;
    data[1616] = -'sd36473;
    data[1617] = -'sd18524;
    data[1618] =  'sd71221;
    data[1619] =  'sd28423;
    data[1620] = -'sd21726;
    data[1621] =  'sd55211;
    data[1622] = -'sd51627;
    data[1623] =  'sd69547;
    data[1624] =  'sd20053;
    data[1625] = -'sd63576;
    data[1626] =  'sd9802;
    data[1627] =  'sd49010;
    data[1628] =  'sd81209;
    data[1629] =  'sd78363;
    data[1630] =  'sd64133;
    data[1631] = -'sd7017;
    data[1632] = -'sd35085;
    data[1633] = -'sd11584;
    data[1634] = -'sd57920;
    data[1635] =  'sd38082;
    data[1636] =  'sd26569;
    data[1637] = -'sd30996;
    data[1638] =  'sd8861;
    data[1639] =  'sd44305;
    data[1640] =  'sd57684;
    data[1641] = -'sd39262;
    data[1642] = -'sd32469;
    data[1643] =  'sd1496;
    data[1644] =  'sd7480;
    data[1645] =  'sd37400;
    data[1646] =  'sd23159;
    data[1647] = -'sd48046;
    data[1648] = -'sd76389;
    data[1649] = -'sd54263;
    data[1650] =  'sd56367;
    data[1651] = -'sd45847;
    data[1652] = -'sd65394;
    data[1653] =  'sd712;
    data[1654] =  'sd3560;
    data[1655] =  'sd17800;
    data[1656] = -'sd74841;
    data[1657] = -'sd46523;
    data[1658] = -'sd68774;
    data[1659] = -'sd16188;
    data[1660] = -'sd80940;
    data[1661] = -'sd77018;
    data[1662] = -'sd57408;
    data[1663] =  'sd40642;
    data[1664] =  'sd39369;
    data[1665] =  'sd33004;
    data[1666] =  'sd1179;
    data[1667] =  'sd5895;
    data[1668] =  'sd29475;
    data[1669] = -'sd16466;
    data[1670] =  'sd81511;
    data[1671] =  'sd79873;
    data[1672] =  'sd71683;
    data[1673] =  'sd30733;
    data[1674] = -'sd10176;
    data[1675] = -'sd50880;
    data[1676] =  'sd73282;
    data[1677] =  'sd38728;
    data[1678] =  'sd29799;
    data[1679] = -'sd14846;
    data[1680] = -'sd74230;
    data[1681] = -'sd43468;
    data[1682] = -'sd53499;
    data[1683] =  'sd60187;
    data[1684] = -'sd26747;
    data[1685] =  'sd30106;
    data[1686] = -'sd13311;
    data[1687] = -'sd66555;
    data[1688] = -'sd5093;
    data[1689] = -'sd25465;
    data[1690] =  'sd36516;
    data[1691] =  'sd18739;
    data[1692] = -'sd70146;
    data[1693] = -'sd23048;
    data[1694] =  'sd48601;
    data[1695] =  'sd79164;
    data[1696] =  'sd68138;
    data[1697] =  'sd13008;
    data[1698] =  'sd65040;
    data[1699] = -'sd2482;
    data[1700] = -'sd12410;
    data[1701] = -'sd62050;
    data[1702] =  'sd17432;
    data[1703] = -'sd76681;
    data[1704] = -'sd55723;
    data[1705] =  'sd49067;
    data[1706] =  'sd81494;
    data[1707] =  'sd79788;
    data[1708] =  'sd71258;
    data[1709] =  'sd28608;
    data[1710] = -'sd20801;
    data[1711] =  'sd59836;
    data[1712] = -'sd28502;
    data[1713] =  'sd21331;
    data[1714] = -'sd57186;
    data[1715] =  'sd41752;
    data[1716] =  'sd44919;
    data[1717] =  'sd60754;
    data[1718] = -'sd23912;
    data[1719] =  'sd44281;
    data[1720] =  'sd57564;
    data[1721] = -'sd39862;
    data[1722] = -'sd35469;
    data[1723] = -'sd13504;
    data[1724] = -'sd67520;
    data[1725] = -'sd9918;
    data[1726] = -'sd49590;
    data[1727] =  'sd79732;
    data[1728] =  'sd70978;
    data[1729] =  'sd27208;
    data[1730] = -'sd27801;
    data[1731] =  'sd24836;
    data[1732] = -'sd39661;
    data[1733] = -'sd34464;
    data[1734] = -'sd8479;
    data[1735] = -'sd42395;
    data[1736] = -'sd48134;
    data[1737] = -'sd76829;
    data[1738] = -'sd56463;
    data[1739] =  'sd45367;
    data[1740] =  'sd62994;
    data[1741] = -'sd12712;
    data[1742] = -'sd63560;
    data[1743] =  'sd9882;
    data[1744] =  'sd49410;
    data[1745] = -'sd80632;
    data[1746] = -'sd75478;
    data[1747] = -'sd49708;
    data[1748] =  'sd79142;
    data[1749] =  'sd68028;
    data[1750] =  'sd12458;
    data[1751] =  'sd62290;
    data[1752] = -'sd16232;
    data[1753] = -'sd81160;
    data[1754] = -'sd78118;
    data[1755] = -'sd62908;
    data[1756] =  'sd13142;
    data[1757] =  'sd65710;
    data[1758] =  'sd868;
    data[1759] =  'sd4340;
    data[1760] =  'sd21700;
    data[1761] = -'sd55341;
    data[1762] =  'sd50977;
    data[1763] = -'sd72797;
    data[1764] = -'sd36303;
    data[1765] = -'sd17674;
    data[1766] =  'sd75471;
    data[1767] =  'sd49673;
    data[1768] = -'sd79317;
    data[1769] = -'sd68903;
    data[1770] = -'sd16833;
    data[1771] =  'sd79676;
    data[1772] =  'sd70698;
    data[1773] =  'sd25808;
    data[1774] = -'sd34801;
    data[1775] = -'sd10164;
    data[1776] = -'sd50820;
    data[1777] =  'sd73582;
    data[1778] =  'sd40228;
    data[1779] =  'sd37299;
    data[1780] =  'sd22654;
    data[1781] = -'sd50571;
    data[1782] =  'sd74827;
    data[1783] =  'sd46453;
    data[1784] =  'sd68424;
    data[1785] =  'sd14438;
    data[1786] =  'sd72190;
    data[1787] =  'sd33268;
    data[1788] =  'sd2499;
    data[1789] =  'sd12495;
    data[1790] =  'sd62475;
    data[1791] = -'sd15307;
    data[1792] = -'sd76535;
    data[1793] = -'sd54993;
    data[1794] =  'sd52717;
    data[1795] = -'sd64097;
    data[1796] =  'sd7197;
    data[1797] =  'sd35985;
    data[1798] =  'sd16084;
    data[1799] =  'sd80420;
    data[1800] =  'sd74418;
    data[1801] =  'sd44408;
    data[1802] =  'sd58199;
    data[1803] = -'sd36687;
    data[1804] = -'sd19594;
    data[1805] =  'sd65871;
    data[1806] =  'sd1673;
    data[1807] =  'sd8365;
    data[1808] =  'sd41825;
    data[1809] =  'sd45284;
    data[1810] =  'sd62579;
    data[1811] = -'sd14787;
    data[1812] = -'sd73935;
    data[1813] = -'sd41993;
    data[1814] = -'sd46124;
    data[1815] = -'sd66779;
    data[1816] = -'sd6213;
    data[1817] = -'sd31065;
    data[1818] =  'sd8516;
    data[1819] =  'sd42580;
    data[1820] =  'sd49059;
    data[1821] =  'sd81454;
    data[1822] =  'sd79588;
    data[1823] =  'sd70258;
    data[1824] =  'sd23608;
    data[1825] = -'sd45801;
    data[1826] = -'sd65164;
    data[1827] =  'sd1862;
    data[1828] =  'sd9310;
    data[1829] =  'sd46550;
    data[1830] =  'sd68909;
    data[1831] =  'sd16863;
    data[1832] = -'sd79526;
    data[1833] = -'sd69948;
    data[1834] = -'sd22058;
    data[1835] =  'sd53551;
    data[1836] = -'sd59927;
    data[1837] =  'sd28047;
    data[1838] = -'sd23606;
    data[1839] =  'sd45811;
    data[1840] =  'sd65214;
    data[1841] = -'sd1612;
    data[1842] = -'sd8060;
    data[1843] = -'sd40300;
    data[1844] = -'sd37659;
    data[1845] = -'sd24454;
    data[1846] =  'sd41571;
    data[1847] =  'sd44014;
    data[1848] =  'sd56229;
    data[1849] = -'sd46537;
    data[1850] = -'sd68844;
    data[1851] = -'sd16538;
    data[1852] =  'sd81151;
    data[1853] =  'sd78073;
    data[1854] =  'sd62683;
    data[1855] = -'sd14267;
    data[1856] = -'sd71335;
    data[1857] = -'sd28993;
    data[1858] =  'sd18876;
    data[1859] = -'sd69461;
    data[1860] = -'sd19623;
    data[1861] =  'sd65726;
    data[1862] =  'sd948;
    data[1863] =  'sd4740;
    data[1864] =  'sd23700;
    data[1865] = -'sd45341;
    data[1866] = -'sd62864;
    data[1867] =  'sd13362;
    data[1868] =  'sd66810;
    data[1869] =  'sd6368;
    data[1870] =  'sd31840;
    data[1871] = -'sd4641;
    data[1872] = -'sd23205;
    data[1873] =  'sd47816;
    data[1874] =  'sd75239;
    data[1875] =  'sd48513;
    data[1876] =  'sd78724;
    data[1877] =  'sd65938;
    data[1878] =  'sd2008;
    data[1879] =  'sd10040;
    data[1880] =  'sd50200;
    data[1881] = -'sd76682;
    data[1882] = -'sd55728;
    data[1883] =  'sd49042;
    data[1884] =  'sd81369;
    data[1885] =  'sd79163;
    data[1886] =  'sd68133;
    data[1887] =  'sd12983;
    data[1888] =  'sd64915;
    data[1889] = -'sd3107;
    data[1890] = -'sd15535;
    data[1891] = -'sd77675;
    data[1892] = -'sd60693;
    data[1893] =  'sd24217;
    data[1894] = -'sd42756;
    data[1895] = -'sd49939;
    data[1896] =  'sd77987;
    data[1897] =  'sd62253;
    data[1898] = -'sd16417;
    data[1899] =  'sd81756;
    data[1900] =  'sd81098;
    data[1901] =  'sd77808;
    data[1902] =  'sd61358;
    data[1903] = -'sd20892;
    data[1904] =  'sd59381;
    data[1905] = -'sd30777;
    data[1906] =  'sd9956;
    data[1907] =  'sd49780;
    data[1908] = -'sd78782;
    data[1909] = -'sd66228;
    data[1910] = -'sd3458;
    data[1911] = -'sd17290;
    data[1912] =  'sd77391;
    data[1913] =  'sd59273;
    data[1914] = -'sd31317;
    data[1915] =  'sd7256;
    data[1916] =  'sd36280;
    data[1917] =  'sd17559;
    data[1918] = -'sd76046;
    data[1919] = -'sd52548;
    data[1920] =  'sd64942;
    data[1921] = -'sd2972;
    data[1922] = -'sd14860;
    data[1923] = -'sd74300;
    data[1924] = -'sd43818;
    data[1925] = -'sd55249;
    data[1926] =  'sd51437;
    data[1927] = -'sd70497;
    data[1928] = -'sd24803;
    data[1929] =  'sd39826;
    data[1930] =  'sd35289;
    data[1931] =  'sd12604;
    data[1932] =  'sd63020;
    data[1933] = -'sd12582;
    data[1934] = -'sd62910;
    data[1935] =  'sd13132;
    data[1936] =  'sd65660;
    data[1937] =  'sd618;
    data[1938] =  'sd3090;
    data[1939] =  'sd15450;
    data[1940] =  'sd77250;
    data[1941] =  'sd58568;
    data[1942] = -'sd34842;
    data[1943] = -'sd10369;
    data[1944] = -'sd51845;
    data[1945] =  'sd68457;
    data[1946] =  'sd14603;
    data[1947] =  'sd73015;
    data[1948] =  'sd37393;
    data[1949] =  'sd23124;
    data[1950] = -'sd48221;
    data[1951] = -'sd77264;
    data[1952] = -'sd58638;
    data[1953] =  'sd34492;
    data[1954] =  'sd8619;
    data[1955] =  'sd43095;
    data[1956] =  'sd51634;
    data[1957] = -'sd69512;
    data[1958] = -'sd19878;
    data[1959] =  'sd64451;
    data[1960] = -'sd5427;
    data[1961] = -'sd27135;
    data[1962] =  'sd28166;
    data[1963] = -'sd23011;
    data[1964] =  'sd48786;
    data[1965] =  'sd80089;
    data[1966] =  'sd72763;
    data[1967] =  'sd36133;
    data[1968] =  'sd16824;
    data[1969] = -'sd79721;
    data[1970] = -'sd70923;
    data[1971] = -'sd26933;
    data[1972] =  'sd29176;
    data[1973] = -'sd17961;
    data[1974] =  'sd74036;
    data[1975] =  'sd42498;
    data[1976] =  'sd48649;
    data[1977] =  'sd79404;
    data[1978] =  'sd69338;
    data[1979] =  'sd19008;
    data[1980] = -'sd68801;
    data[1981] = -'sd16323;
    data[1982] = -'sd81615;
    data[1983] = -'sd80393;
    data[1984] = -'sd74283;
    data[1985] = -'sd43733;
    data[1986] = -'sd54824;
    data[1987] =  'sd53562;
    data[1988] = -'sd59872;
    data[1989] =  'sd28322;
    data[1990] = -'sd22231;
    data[1991] =  'sd52686;
    data[1992] = -'sd64252;
    data[1993] =  'sd6422;
    data[1994] =  'sd32110;
    data[1995] = -'sd3291;
    data[1996] = -'sd16455;
    data[1997] =  'sd81566;
    data[1998] =  'sd80148;
    data[1999] =  'sd73058;
    data[2000] =  'sd37608;
    data[2001] =  'sd24199;
    data[2002] = -'sd42846;
    data[2003] = -'sd50389;
    data[2004] =  'sd75737;
    data[2005] =  'sd51003;
    data[2006] = -'sd72667;
    data[2007] = -'sd35653;
    data[2008] = -'sd14424;
    data[2009] = -'sd72120;
    data[2010] = -'sd32918;
    data[2011] = -'sd749;
    data[2012] = -'sd3745;
    data[2013] = -'sd18725;
    data[2014] =  'sd70216;
    data[2015] =  'sd23398;
    data[2016] = -'sd46851;
    data[2017] = -'sd70414;
    data[2018] = -'sd24388;
    data[2019] =  'sd41901;
    data[2020] =  'sd45664;
    data[2021] =  'sd64479;
    data[2022] = -'sd5287;
    data[2023] = -'sd26435;
    data[2024] =  'sd31666;
    data[2025] = -'sd5511;
    data[2026] = -'sd27555;
    data[2027] =  'sd26066;
    data[2028] = -'sd33511;
    data[2029] = -'sd3714;
    data[2030] = -'sd18570;
    data[2031] =  'sd70991;
    data[2032] =  'sd27273;
    data[2033] = -'sd27476;
    data[2034] =  'sd26461;
    data[2035] = -'sd31536;
    data[2036] =  'sd6161;
    data[2037] =  'sd30805;
    data[2038] = -'sd9816;
    data[2039] = -'sd49080;
    data[2040] = -'sd81559;
    data[2041] = -'sd80113;
    data[2042] = -'sd72883;
    data[2043] = -'sd36733;
    data[2044] = -'sd19824;
    data[2045] =  'sd64721;
    data[2046] = -'sd4077;
    data[2047] = -'sd20385;
    data[2048] =  'sd61916;
    data[2049] = -'sd18102;
    data[2050] =  'sd73331;
    data[2051] =  'sd38973;
    data[2052] =  'sd31024;
    data[2053] = -'sd8721;
    data[2054] = -'sd43605;
    data[2055] = -'sd54184;
    data[2056] =  'sd56762;
    data[2057] = -'sd43872;
    data[2058] = -'sd55519;
    data[2059] =  'sd50087;
    data[2060] = -'sd77247;
    data[2061] = -'sd58553;
    data[2062] =  'sd34917;
    data[2063] =  'sd10744;
    data[2064] =  'sd53720;
    data[2065] = -'sd59082;
    data[2066] =  'sd32272;
    data[2067] = -'sd2481;
    data[2068] = -'sd12405;
    data[2069] = -'sd62025;
    data[2070] =  'sd17557;
    data[2071] = -'sd76056;
    data[2072] = -'sd52598;
    data[2073] =  'sd64692;
    data[2074] = -'sd4222;
    data[2075] = -'sd21110;
    data[2076] =  'sd58291;
    data[2077] = -'sd36227;
    data[2078] = -'sd17294;
    data[2079] =  'sd77371;
    data[2080] =  'sd59173;
    data[2081] = -'sd31817;
    data[2082] =  'sd4756;
    data[2083] =  'sd23780;
    data[2084] = -'sd44941;
    data[2085] = -'sd60864;
    data[2086] =  'sd23362;
    data[2087] = -'sd47031;
    data[2088] = -'sd71314;
    data[2089] = -'sd28888;
    data[2090] =  'sd19401;
    data[2091] = -'sd66836;
    data[2092] = -'sd6498;
    data[2093] = -'sd32490;
    data[2094] =  'sd1391;
    data[2095] =  'sd6955;
    data[2096] =  'sd34775;
    data[2097] =  'sd10034;
    data[2098] =  'sd50170;
    data[2099] = -'sd76832;
    data[2100] = -'sd56478;
    data[2101] =  'sd45292;
    data[2102] =  'sd62619;
    data[2103] = -'sd14587;
    data[2104] = -'sd72935;
    data[2105] = -'sd36993;
    data[2106] = -'sd21124;
    data[2107] =  'sd58221;
    data[2108] = -'sd36577;
    data[2109] = -'sd19044;
    data[2110] =  'sd68621;
    data[2111] =  'sd15423;
    data[2112] =  'sd77115;
    data[2113] =  'sd57893;
    data[2114] = -'sd38217;
    data[2115] = -'sd27244;
    data[2116] =  'sd27621;
    data[2117] = -'sd25736;
    data[2118] =  'sd35161;
    data[2119] =  'sd11964;
    data[2120] =  'sd59820;
    data[2121] = -'sd28582;
    data[2122] =  'sd20931;
    data[2123] = -'sd59186;
    data[2124] =  'sd31752;
    data[2125] = -'sd5081;
    data[2126] = -'sd25405;
    data[2127] =  'sd36816;
    data[2128] =  'sd20239;
    data[2129] = -'sd62646;
    data[2130] =  'sd14452;
    data[2131] =  'sd72260;
    data[2132] =  'sd33618;
    data[2133] =  'sd4249;
    data[2134] =  'sd21245;
    data[2135] = -'sd57616;
    data[2136] =  'sd39602;
    data[2137] =  'sd34169;
    data[2138] =  'sd7004;
    data[2139] =  'sd35020;
    data[2140] =  'sd11259;
    data[2141] =  'sd56295;
    data[2142] = -'sd46207;
    data[2143] = -'sd67194;
    data[2144] = -'sd8288;
    data[2145] = -'sd41440;
    data[2146] = -'sd43359;
    data[2147] = -'sd52954;
    data[2148] =  'sd62912;
    data[2149] = -'sd13122;
    data[2150] = -'sd65610;
    data[2151] = -'sd368;
    data[2152] = -'sd1840;
    data[2153] = -'sd9200;
    data[2154] = -'sd46000;
    data[2155] = -'sd66159;
    data[2156] = -'sd3113;
    data[2157] = -'sd15565;
    data[2158] = -'sd77825;
    data[2159] = -'sd61443;
    data[2160] =  'sd20467;
    data[2161] = -'sd61506;
    data[2162] =  'sd20152;
    data[2163] = -'sd63081;
    data[2164] =  'sd12277;
    data[2165] =  'sd61385;
    data[2166] = -'sd20757;
    data[2167] =  'sd60056;
    data[2168] = -'sd27402;
    data[2169] =  'sd26831;
    data[2170] = -'sd29686;
    data[2171] =  'sd15411;
    data[2172] =  'sd77055;
    data[2173] =  'sd57593;
    data[2174] = -'sd39717;
    data[2175] = -'sd34744;
    data[2176] = -'sd9879;
    data[2177] = -'sd49395;
    data[2178] =  'sd80707;
    data[2179] =  'sd75853;
    data[2180] =  'sd51583;
    data[2181] = -'sd69767;
    data[2182] = -'sd21153;
    data[2183] =  'sd58076;
    data[2184] = -'sd37302;
    data[2185] = -'sd22669;
    data[2186] =  'sd50496;
    data[2187] = -'sd75202;
    data[2188] = -'sd48328;
    data[2189] = -'sd77799;
    data[2190] = -'sd61313;
    data[2191] =  'sd21117;
    data[2192] = -'sd58256;
    data[2193] =  'sd36402;
    data[2194] =  'sd18169;
    data[2195] = -'sd72996;
    data[2196] = -'sd37298;
    data[2197] = -'sd22649;
    data[2198] =  'sd50596;
    data[2199] = -'sd74702;
    data[2200] = -'sd45828;
    data[2201] = -'sd65299;
    data[2202] =  'sd1187;
    data[2203] =  'sd5935;
    data[2204] =  'sd29675;
    data[2205] = -'sd15466;
    data[2206] = -'sd77330;
    data[2207] = -'sd58968;
    data[2208] =  'sd32842;
    data[2209] =  'sd369;
    data[2210] =  'sd1845;
    data[2211] =  'sd9225;
    data[2212] =  'sd46125;
    data[2213] =  'sd66784;
    data[2214] =  'sd6238;
    data[2215] =  'sd31190;
    data[2216] = -'sd7891;
    data[2217] = -'sd39455;
    data[2218] = -'sd33434;
    data[2219] = -'sd3329;
    data[2220] = -'sd16645;
    data[2221] =  'sd80616;
    data[2222] =  'sd75398;
    data[2223] =  'sd49308;
    data[2224] = -'sd81142;
    data[2225] = -'sd78028;
    data[2226] = -'sd62458;
    data[2227] =  'sd15392;
    data[2228] =  'sd76960;
    data[2229] =  'sd57118;
    data[2230] = -'sd42092;
    data[2231] = -'sd46619;
    data[2232] = -'sd69254;
    data[2233] = -'sd18588;
    data[2234] =  'sd70901;
    data[2235] =  'sd26823;
    data[2236] = -'sd29726;
    data[2237] =  'sd15211;
    data[2238] =  'sd76055;
    data[2239] =  'sd52593;
    data[2240] = -'sd64717;
    data[2241] =  'sd4097;
    data[2242] =  'sd20485;
    data[2243] = -'sd61416;
    data[2244] =  'sd20602;
    data[2245] = -'sd60831;
    data[2246] =  'sd23527;
    data[2247] = -'sd46206;
    data[2248] = -'sd67189;
    data[2249] = -'sd8263;
    data[2250] = -'sd41315;
    data[2251] = -'sd42734;
    data[2252] = -'sd49829;
    data[2253] =  'sd78537;
    data[2254] =  'sd65003;
    data[2255] = -'sd2667;
    data[2256] = -'sd13335;
    data[2257] = -'sd66675;
    data[2258] = -'sd5693;
    data[2259] = -'sd28465;
    data[2260] =  'sd21516;
    data[2261] = -'sd56261;
    data[2262] =  'sd46377;
    data[2263] =  'sd68044;
    data[2264] =  'sd12538;
    data[2265] =  'sd62690;
    data[2266] = -'sd14232;
    data[2267] = -'sd71160;
    data[2268] = -'sd28118;
    data[2269] =  'sd23251;
    data[2270] = -'sd47586;
    data[2271] = -'sd74089;
    data[2272] = -'sd42763;
    data[2273] = -'sd49974;
    data[2274] =  'sd77812;
    data[2275] =  'sd61378;
    data[2276] = -'sd20792;
    data[2277] =  'sd59881;
    data[2278] = -'sd28277;
    data[2279] =  'sd22456;
    data[2280] = -'sd51561;
    data[2281] =  'sd69877;
    data[2282] =  'sd21703;
    data[2283] = -'sd55326;
    data[2284] =  'sd51052;
    data[2285] = -'sd72422;
    data[2286] = -'sd34428;
    data[2287] = -'sd8299;
    data[2288] = -'sd41495;
    data[2289] = -'sd43634;
    data[2290] = -'sd54329;
    data[2291] =  'sd56037;
    data[2292] = -'sd47497;
    data[2293] = -'sd73644;
    data[2294] = -'sd40538;
    data[2295] = -'sd38849;
    data[2296] = -'sd30404;
    data[2297] =  'sd11821;
    data[2298] =  'sd59105;
    data[2299] = -'sd32157;
    data[2300] =  'sd3056;
    data[2301] =  'sd15280;
    data[2302] =  'sd76400;
    data[2303] =  'sd54318;
    data[2304] = -'sd56092;
    data[2305] =  'sd47222;
    data[2306] =  'sd72269;
    data[2307] =  'sd33663;
    data[2308] =  'sd4474;
    data[2309] =  'sd22370;
    data[2310] = -'sd51991;
    data[2311] =  'sd67727;
    data[2312] =  'sd10953;
    data[2313] =  'sd54765;
    data[2314] = -'sd53857;
    data[2315] =  'sd58397;
    data[2316] = -'sd35697;
    data[2317] = -'sd14644;
    data[2318] = -'sd73220;
    data[2319] = -'sd38418;
    data[2320] = -'sd28249;
    data[2321] =  'sd22596;
    data[2322] = -'sd50861;
    data[2323] =  'sd73377;
    data[2324] =  'sd39203;
    data[2325] =  'sd32174;
    data[2326] = -'sd2971;
    data[2327] = -'sd14855;
    data[2328] = -'sd74275;
    data[2329] = -'sd43693;
    data[2330] = -'sd54624;
    data[2331] =  'sd54562;
    data[2332] = -'sd54872;
    data[2333] =  'sd53322;
    data[2334] = -'sd61072;
    data[2335] =  'sd22322;
    data[2336] = -'sd52231;
    data[2337] =  'sd66527;
    data[2338] =  'sd4953;
    data[2339] =  'sd24765;
    data[2340] = -'sd40016;
    data[2341] = -'sd36239;
    data[2342] = -'sd17354;
    data[2343] =  'sd77071;
    data[2344] =  'sd57673;
    data[2345] = -'sd39317;
    data[2346] = -'sd32744;
    data[2347] =  'sd121;
    data[2348] =  'sd605;
    data[2349] =  'sd3025;
    data[2350] =  'sd15125;
    data[2351] =  'sd75625;
    data[2352] =  'sd50443;
    data[2353] = -'sd75467;
    data[2354] = -'sd49653;
    data[2355] =  'sd79417;
    data[2356] =  'sd69403;
    data[2357] =  'sd19333;
    data[2358] = -'sd67176;
    data[2359] = -'sd8198;
    data[2360] = -'sd40990;
    data[2361] = -'sd41109;
    data[2362] = -'sd41704;
    data[2363] = -'sd44679;
    data[2364] = -'sd59554;
    data[2365] =  'sd29912;
    data[2366] = -'sd14281;
    data[2367] = -'sd71405;
    data[2368] = -'sd29343;
    data[2369] =  'sd17126;
    data[2370] = -'sd78211;
    data[2371] = -'sd63373;
    data[2372] =  'sd10817;
    data[2373] =  'sd54085;
    data[2374] = -'sd57257;
    data[2375] =  'sd41397;
    data[2376] =  'sd43144;
    data[2377] =  'sd51879;
    data[2378] = -'sd68287;
    data[2379] = -'sd13753;
    data[2380] = -'sd68765;
    data[2381] = -'sd16143;
    data[2382] = -'sd80715;
    data[2383] = -'sd75893;
    data[2384] = -'sd51783;
    data[2385] =  'sd68767;
    data[2386] =  'sd16153;
    data[2387] =  'sd80765;
    data[2388] =  'sd76143;
    data[2389] =  'sd53033;
    data[2390] = -'sd62517;
    data[2391] =  'sd15097;
    data[2392] =  'sd75485;
    data[2393] =  'sd49743;
    data[2394] = -'sd78967;
    data[2395] = -'sd67153;
    data[2396] = -'sd8083;
    data[2397] = -'sd40415;
    data[2398] = -'sd38234;
    data[2399] = -'sd27329;
    data[2400] =  'sd27196;
    data[2401] = -'sd27861;
    data[2402] =  'sd24536;
    data[2403] = -'sd41161;
    data[2404] = -'sd41964;
    data[2405] = -'sd45979;
    data[2406] = -'sd66054;
    data[2407] = -'sd2588;
    data[2408] = -'sd12940;
    data[2409] = -'sd64700;
    data[2410] =  'sd4182;
    data[2411] =  'sd20910;
    data[2412] = -'sd59291;
    data[2413] =  'sd31227;
    data[2414] = -'sd7706;
    data[2415] = -'sd38530;
    data[2416] = -'sd28809;
    data[2417] =  'sd19796;
    data[2418] = -'sd64861;
    data[2419] =  'sd3377;
    data[2420] =  'sd16885;
    data[2421] = -'sd79416;
    data[2422] = -'sd69398;
    data[2423] = -'sd19308;
    data[2424] =  'sd67301;
    data[2425] =  'sd8823;
    data[2426] =  'sd44115;
    data[2427] =  'sd56734;
    data[2428] = -'sd44012;
    data[2429] = -'sd56219;
    data[2430] =  'sd46587;
    data[2431] =  'sd69094;
    data[2432] =  'sd17788;
    data[2433] = -'sd74901;
    data[2434] = -'sd46823;
    data[2435] = -'sd70274;
    data[2436] = -'sd23688;
    data[2437] =  'sd45401;
    data[2438] =  'sd63164;
    data[2439] = -'sd11862;
    data[2440] = -'sd59310;
    data[2441] =  'sd31132;
    data[2442] = -'sd8181;
    data[2443] = -'sd40905;
    data[2444] = -'sd40684;
    data[2445] = -'sd39579;
    data[2446] = -'sd34054;
    data[2447] = -'sd6429;
    data[2448] = -'sd32145;
    data[2449] =  'sd3116;
    data[2450] =  'sd15580;
    data[2451] =  'sd77900;
    data[2452] =  'sd61818;
    data[2453] = -'sd18592;
    data[2454] =  'sd70881;
    data[2455] =  'sd26723;
    data[2456] = -'sd30226;
    data[2457] =  'sd12711;
    data[2458] =  'sd63555;
    data[2459] = -'sd9907;
    data[2460] = -'sd49535;
    data[2461] =  'sd80007;
    data[2462] =  'sd72353;
    data[2463] =  'sd34083;
    data[2464] =  'sd6574;
    data[2465] =  'sd32870;
    data[2466] =  'sd509;
    data[2467] =  'sd2545;
    data[2468] =  'sd12725;
    data[2469] =  'sd63625;
    data[2470] = -'sd9557;
    data[2471] = -'sd47785;
    data[2472] = -'sd75084;
    data[2473] = -'sd47738;
    data[2474] = -'sd74849;
    data[2475] = -'sd46563;
    data[2476] = -'sd68974;
    data[2477] = -'sd17188;
    data[2478] =  'sd77901;
    data[2479] =  'sd61823;
    data[2480] = -'sd18567;
    data[2481] =  'sd71006;
    data[2482] =  'sd27348;
    data[2483] = -'sd27101;
    data[2484] =  'sd28336;
    data[2485] = -'sd22161;
    data[2486] =  'sd53036;
    data[2487] = -'sd62502;
    data[2488] =  'sd15172;
    data[2489] =  'sd75860;
    data[2490] =  'sd51618;
    data[2491] = -'sd69592;
    data[2492] = -'sd20278;
    data[2493] =  'sd62451;
    data[2494] = -'sd15427;
    data[2495] = -'sd77135;
    data[2496] = -'sd57993;
    data[2497] =  'sd37717;
    data[2498] =  'sd24744;
    data[2499] = -'sd40121;
    data[2500] = -'sd36764;
    data[2501] = -'sd19979;
    data[2502] =  'sd63946;
    data[2503] = -'sd7952;
    data[2504] = -'sd39760;
    data[2505] = -'sd34959;
    data[2506] = -'sd10954;
    data[2507] = -'sd54770;
    data[2508] =  'sd53832;
    data[2509] = -'sd58522;
    data[2510] =  'sd35072;
    data[2511] =  'sd11519;
    data[2512] =  'sd57595;
    data[2513] = -'sd39707;
    data[2514] = -'sd34694;
    data[2515] = -'sd9629;
    data[2516] = -'sd48145;
    data[2517] = -'sd76884;
    data[2518] = -'sd56738;
    data[2519] =  'sd43992;
    data[2520] =  'sd56119;
    data[2521] = -'sd47087;
    data[2522] = -'sd71594;
    data[2523] = -'sd30288;
    data[2524] =  'sd12401;
    data[2525] =  'sd62005;
    data[2526] = -'sd17657;
    data[2527] =  'sd75556;
    data[2528] =  'sd50098;
    data[2529] = -'sd77192;
    data[2530] = -'sd58278;
    data[2531] =  'sd36292;
    data[2532] =  'sd17619;
    data[2533] = -'sd75746;
    data[2534] = -'sd51048;
    data[2535] =  'sd72442;
    data[2536] =  'sd34528;
    data[2537] =  'sd8799;
    data[2538] =  'sd43995;
    data[2539] =  'sd56134;
    data[2540] = -'sd47012;
    data[2541] = -'sd71219;
    data[2542] = -'sd28413;
    data[2543] =  'sd21776;
    data[2544] = -'sd54961;
    data[2545] =  'sd52877;
    data[2546] = -'sd63297;
    data[2547] =  'sd11197;
    data[2548] =  'sd55985;
    data[2549] = -'sd47757;
    data[2550] = -'sd74944;
    data[2551] = -'sd47038;
    data[2552] = -'sd71349;
    data[2553] = -'sd29063;
    data[2554] =  'sd18526;
    data[2555] = -'sd71211;
    data[2556] = -'sd28373;
    data[2557] =  'sd21976;
    data[2558] = -'sd53961;
    data[2559] =  'sd57877;
    data[2560] = -'sd38297;
    data[2561] = -'sd27644;
    data[2562] =  'sd25621;
    data[2563] = -'sd35736;
    data[2564] = -'sd14839;
    data[2565] = -'sd74195;
    data[2566] = -'sd43293;
    data[2567] = -'sd52624;
    data[2568] =  'sd64562;
    data[2569] = -'sd4872;
    data[2570] = -'sd24360;
    data[2571] =  'sd42041;
    data[2572] =  'sd46364;
    data[2573] =  'sd67979;
    data[2574] =  'sd12213;
    data[2575] =  'sd61065;
    data[2576] = -'sd22357;
    data[2577] =  'sd52056;
    data[2578] = -'sd67402;
    data[2579] = -'sd9328;
    data[2580] = -'sd46640;
    data[2581] = -'sd69359;
    data[2582] = -'sd19113;
    data[2583] =  'sd68276;
    data[2584] =  'sd13698;
    data[2585] =  'sd68490;
    data[2586] =  'sd14768;
    data[2587] =  'sd73840;
    data[2588] =  'sd41518;
    data[2589] =  'sd43749;
    data[2590] =  'sd54904;
    data[2591] = -'sd53162;
    data[2592] =  'sd61872;
    data[2593] = -'sd18322;
    data[2594] =  'sd72231;
    data[2595] =  'sd33473;
    data[2596] =  'sd3524;
    data[2597] =  'sd17620;
    data[2598] = -'sd75741;
    data[2599] = -'sd51023;
    data[2600] =  'sd72567;
    data[2601] =  'sd35153;
    data[2602] =  'sd11924;
    data[2603] =  'sd59620;
    data[2604] = -'sd29582;
    data[2605] =  'sd15931;
    data[2606] =  'sd79655;
    data[2607] =  'sd70593;
    data[2608] =  'sd25283;
    data[2609] = -'sd37426;
    data[2610] = -'sd23289;
    data[2611] =  'sd47396;
    data[2612] =  'sd73139;
    data[2613] =  'sd38013;
    data[2614] =  'sd26224;
    data[2615] = -'sd32721;
    data[2616] =  'sd236;
    data[2617] =  'sd1180;
    data[2618] =  'sd5900;
    data[2619] =  'sd29500;
    data[2620] = -'sd16341;
    data[2621] = -'sd81705;
    data[2622] = -'sd80843;
    data[2623] = -'sd76533;
    data[2624] = -'sd54983;
    data[2625] =  'sd52767;
    data[2626] = -'sd63847;
    data[2627] =  'sd8447;
    data[2628] =  'sd42235;
    data[2629] =  'sd47334;
    data[2630] =  'sd72829;
    data[2631] =  'sd36463;
    data[2632] =  'sd18474;
    data[2633] = -'sd71471;
    data[2634] = -'sd29673;
    data[2635] =  'sd15476;
    data[2636] =  'sd77380;
    data[2637] =  'sd59218;
    data[2638] = -'sd31592;
    data[2639] =  'sd5881;
    data[2640] =  'sd29405;
    data[2641] = -'sd16816;
    data[2642] =  'sd79761;
    data[2643] =  'sd71123;
    data[2644] =  'sd27933;
    data[2645] = -'sd24176;
    data[2646] =  'sd42961;
    data[2647] =  'sd50964;
    data[2648] = -'sd72862;
    data[2649] = -'sd36628;
    data[2650] = -'sd19299;
    data[2651] =  'sd67346;
    data[2652] =  'sd9048;
    data[2653] =  'sd45240;
    data[2654] =  'sd62359;
    data[2655] = -'sd15887;
    data[2656] = -'sd79435;
    data[2657] = -'sd69493;
    data[2658] = -'sd19783;
    data[2659] =  'sd64926;
    data[2660] = -'sd3052;
    data[2661] = -'sd15260;
    data[2662] = -'sd76300;
    data[2663] = -'sd53818;
    data[2664] =  'sd58592;
    data[2665] = -'sd34722;
    data[2666] = -'sd9769;
    data[2667] = -'sd48845;
    data[2668] = -'sd80384;
    data[2669] = -'sd74238;
    data[2670] = -'sd43508;
    data[2671] = -'sd53699;
    data[2672] =  'sd59187;
    data[2673] = -'sd31747;
    data[2674] =  'sd5106;
    data[2675] =  'sd25530;
    data[2676] = -'sd36191;
    data[2677] = -'sd17114;
    data[2678] =  'sd78271;
    data[2679] =  'sd63673;
    data[2680] = -'sd9317;
    data[2681] = -'sd46585;
    data[2682] = -'sd69084;
    data[2683] = -'sd17738;
    data[2684] =  'sd75151;
    data[2685] =  'sd48073;
    data[2686] =  'sd76524;
    data[2687] =  'sd54938;
    data[2688] = -'sd52992;
    data[2689] =  'sd62722;
    data[2690] = -'sd14072;
    data[2691] = -'sd70360;
    data[2692] = -'sd24118;
    data[2693] =  'sd43251;
    data[2694] =  'sd52414;
    data[2695] = -'sd65612;
    data[2696] = -'sd378;
    data[2697] = -'sd1890;
    data[2698] = -'sd9450;
    data[2699] = -'sd47250;
    data[2700] = -'sd72409;
    data[2701] = -'sd34363;
    data[2702] = -'sd7974;
    data[2703] = -'sd39870;
    data[2704] = -'sd35509;
    data[2705] = -'sd13704;
    data[2706] = -'sd68520;
    data[2707] = -'sd14918;
    data[2708] = -'sd74590;
    data[2709] = -'sd45268;
    data[2710] = -'sd62499;
    data[2711] =  'sd15187;
    data[2712] =  'sd75935;
    data[2713] =  'sd51993;
    data[2714] = -'sd67717;
    data[2715] = -'sd10903;
    data[2716] = -'sd54515;
    data[2717] =  'sd55107;
    data[2718] = -'sd52147;
    data[2719] =  'sd66947;
    data[2720] =  'sd7053;
    data[2721] =  'sd35265;
    data[2722] =  'sd12484;
    data[2723] =  'sd62420;
    data[2724] = -'sd15582;
    data[2725] = -'sd77910;
    data[2726] = -'sd61868;
    data[2727] =  'sd18342;
    data[2728] = -'sd72131;
    data[2729] = -'sd32973;
    data[2730] = -'sd1024;
    data[2731] = -'sd5120;
    data[2732] = -'sd25600;
    data[2733] =  'sd35841;
    data[2734] =  'sd15364;
    data[2735] =  'sd76820;
    data[2736] =  'sd56418;
    data[2737] = -'sd45592;
    data[2738] = -'sd64119;
    data[2739] =  'sd7087;
    data[2740] =  'sd35435;
    data[2741] =  'sd13334;
    data[2742] =  'sd66670;
    data[2743] =  'sd5668;
    data[2744] =  'sd28340;
    data[2745] = -'sd22141;
    data[2746] =  'sd53136;
    data[2747] = -'sd62002;
    data[2748] =  'sd17672;
    data[2749] = -'sd75481;
    data[2750] = -'sd49723;
    data[2751] =  'sd79067;
    data[2752] =  'sd67653;
    data[2753] =  'sd10583;
    data[2754] =  'sd52915;
    data[2755] = -'sd63107;
    data[2756] =  'sd12147;
    data[2757] =  'sd60735;
    data[2758] = -'sd24007;
    data[2759] =  'sd43806;
    data[2760] =  'sd55189;
    data[2761] = -'sd51737;
    data[2762] =  'sd68997;
    data[2763] =  'sd17303;
    data[2764] = -'sd77326;
    data[2765] = -'sd58948;
    data[2766] =  'sd32942;
    data[2767] =  'sd869;
    data[2768] =  'sd4345;
    data[2769] =  'sd21725;
    data[2770] = -'sd55216;
    data[2771] =  'sd51602;
    data[2772] = -'sd69672;
    data[2773] = -'sd20678;
    data[2774] =  'sd60451;
    data[2775] = -'sd25427;
    data[2776] =  'sd36706;
    data[2777] =  'sd19689;
    data[2778] = -'sd65396;
    data[2779] =  'sd702;
    data[2780] =  'sd3510;
    data[2781] =  'sd17550;
    data[2782] = -'sd76091;
    data[2783] = -'sd52773;
    data[2784] =  'sd63817;
    data[2785] = -'sd8597;
    data[2786] = -'sd42985;
    data[2787] = -'sd51084;
    data[2788] =  'sd72262;
    data[2789] =  'sd33628;
    data[2790] =  'sd4299;
    data[2791] =  'sd21495;
    data[2792] = -'sd56366;
    data[2793] =  'sd45852;
    data[2794] =  'sd65419;
    data[2795] = -'sd587;
    data[2796] = -'sd2935;
    data[2797] = -'sd14675;
    data[2798] = -'sd73375;
    data[2799] = -'sd39193;
    data[2800] = -'sd32124;
    data[2801] =  'sd3221;
    data[2802] =  'sd16105;
    data[2803] =  'sd80525;
    data[2804] =  'sd74943;
    data[2805] =  'sd47033;
    data[2806] =  'sd71324;
    data[2807] =  'sd28938;
    data[2808] = -'sd19151;
    data[2809] =  'sd68086;
    data[2810] =  'sd12748;
    data[2811] =  'sd63740;
    data[2812] = -'sd8982;
    data[2813] = -'sd44910;
    data[2814] = -'sd60709;
    data[2815] =  'sd24137;
    data[2816] = -'sd43156;
    data[2817] = -'sd51939;
    data[2818] =  'sd67987;
    data[2819] =  'sd12253;
    data[2820] =  'sd61265;
    data[2821] = -'sd21357;
    data[2822] =  'sd57056;
    data[2823] = -'sd42402;
    data[2824] = -'sd48169;
    data[2825] = -'sd77004;
    data[2826] = -'sd57338;
    data[2827] =  'sd40992;
    data[2828] =  'sd41119;
    data[2829] =  'sd41754;
    data[2830] =  'sd44929;
    data[2831] =  'sd60804;
    data[2832] = -'sd23662;
    data[2833] =  'sd45531;
    data[2834] =  'sd63814;
    data[2835] = -'sd8612;
    data[2836] = -'sd43060;
    data[2837] = -'sd51459;
    data[2838] =  'sd70387;
    data[2839] =  'sd24253;
    data[2840] = -'sd42576;
    data[2841] = -'sd49039;
    data[2842] = -'sd81354;
    data[2843] = -'sd79088;
    data[2844] = -'sd67758;
    data[2845] = -'sd11108;
    data[2846] = -'sd55540;
    data[2847] =  'sd49982;
    data[2848] = -'sd77772;
    data[2849] = -'sd61178;
    data[2850] =  'sd21792;
    data[2851] = -'sd54881;
    data[2852] =  'sd53277;
    data[2853] = -'sd61297;
    data[2854] =  'sd21197;
    data[2855] = -'sd57856;
    data[2856] =  'sd38402;
    data[2857] =  'sd28169;
    data[2858] = -'sd22996;
    data[2859] =  'sd48861;
    data[2860] =  'sd80464;
    data[2861] =  'sd74638;
    data[2862] =  'sd45508;
    data[2863] =  'sd63699;
    data[2864] = -'sd9187;
    data[2865] = -'sd45935;
    data[2866] = -'sd65834;
    data[2867] = -'sd1488;
    data[2868] = -'sd7440;
    data[2869] = -'sd37200;
    data[2870] = -'sd22159;
    data[2871] =  'sd53046;
    data[2872] = -'sd62452;
    data[2873] =  'sd15422;
    data[2874] =  'sd77110;
    data[2875] =  'sd57868;
    data[2876] = -'sd38342;
    data[2877] = -'sd27869;
    data[2878] =  'sd24496;
    data[2879] = -'sd41361;
    data[2880] = -'sd42964;
    data[2881] = -'sd50979;
    data[2882] =  'sd72787;
    data[2883] =  'sd36253;
    data[2884] =  'sd17424;
    data[2885] = -'sd76721;
    data[2886] = -'sd55923;
    data[2887] =  'sd48067;
    data[2888] =  'sd76494;
    data[2889] =  'sd54788;
    data[2890] = -'sd53742;
    data[2891] =  'sd58972;
    data[2892] = -'sd32822;
    data[2893] = -'sd269;
    data[2894] = -'sd1345;
    data[2895] = -'sd6725;
    data[2896] = -'sd33625;
    data[2897] = -'sd4284;
    data[2898] = -'sd21420;
    data[2899] =  'sd56741;
    data[2900] = -'sd43977;
    data[2901] = -'sd56044;
    data[2902] =  'sd47462;
    data[2903] =  'sd73469;
    data[2904] =  'sd39663;
    data[2905] =  'sd34474;
    data[2906] =  'sd8529;
    data[2907] =  'sd42645;
    data[2908] =  'sd49384;
    data[2909] = -'sd80762;
    data[2910] = -'sd76128;
    data[2911] = -'sd52958;
    data[2912] =  'sd62892;
    data[2913] = -'sd13222;
    data[2914] = -'sd66110;
    data[2915] = -'sd2868;
    data[2916] = -'sd14340;
    data[2917] = -'sd71700;
    data[2918] = -'sd30818;
    data[2919] =  'sd9751;
    data[2920] =  'sd48755;
    data[2921] =  'sd79934;
    data[2922] =  'sd71988;
    data[2923] =  'sd32258;
    data[2924] = -'sd2551;
    data[2925] = -'sd12755;
    data[2926] = -'sd63775;
    data[2927] =  'sd8807;
    data[2928] =  'sd44035;
    data[2929] =  'sd56334;
    data[2930] = -'sd46012;
    data[2931] = -'sd66219;
    data[2932] = -'sd3413;
    data[2933] = -'sd17065;
    data[2934] =  'sd78516;
    data[2935] =  'sd64898;
    data[2936] = -'sd3192;
    data[2937] = -'sd15960;
    data[2938] = -'sd79800;
    data[2939] = -'sd71318;
    data[2940] = -'sd28908;
    data[2941] =  'sd19301;
    data[2942] = -'sd67336;
    data[2943] = -'sd8998;
    data[2944] = -'sd44990;
    data[2945] = -'sd61109;
    data[2946] =  'sd22137;
    data[2947] = -'sd53156;
    data[2948] =  'sd61902;
    data[2949] = -'sd18172;
    data[2950] =  'sd72981;
    data[2951] =  'sd37223;
    data[2952] =  'sd22274;
    data[2953] = -'sd52471;
    data[2954] =  'sd65327;
    data[2955] = -'sd1047;
    data[2956] = -'sd5235;
    data[2957] = -'sd26175;
    data[2958] =  'sd32966;
    data[2959] =  'sd989;
    data[2960] =  'sd4945;
    data[2961] =  'sd24725;
    data[2962] = -'sd40216;
    data[2963] = -'sd37239;
    data[2964] = -'sd22354;
    data[2965] =  'sd52071;
    data[2966] = -'sd67327;
    data[2967] = -'sd8953;
    data[2968] = -'sd44765;
    data[2969] = -'sd59984;
    data[2970] =  'sd27762;
    data[2971] = -'sd25031;
    data[2972] =  'sd38686;
    data[2973] =  'sd29589;
    data[2974] = -'sd15896;
    data[2975] = -'sd79480;
    data[2976] = -'sd69718;
    data[2977] = -'sd20908;
    data[2978] =  'sd59301;
    data[2979] = -'sd31177;
    data[2980] =  'sd7956;
    data[2981] =  'sd39780;
    data[2982] =  'sd35059;
    data[2983] =  'sd11454;
    data[2984] =  'sd57270;
    data[2985] = -'sd41332;
    data[2986] = -'sd42819;
    data[2987] = -'sd50254;
    data[2988] =  'sd76412;
    data[2989] =  'sd54378;
    data[2990] = -'sd55792;
    data[2991] =  'sd48722;
    data[2992] =  'sd79769;
    data[2993] =  'sd71163;
    data[2994] =  'sd28133;
    data[2995] = -'sd23176;
    data[2996] =  'sd47961;
    data[2997] =  'sd75964;
    data[2998] =  'sd52138;
    data[2999] = -'sd66992;
    data[3000] = -'sd7278;
    data[3001] = -'sd36390;
    data[3002] = -'sd18109;
    data[3003] =  'sd73296;
    data[3004] =  'sd38798;
    data[3005] =  'sd30149;
    data[3006] = -'sd13096;
    data[3007] = -'sd65480;
    data[3008] =  'sd282;
    data[3009] =  'sd1410;
    data[3010] =  'sd7050;
    data[3011] =  'sd35250;
    data[3012] =  'sd12409;
    data[3013] =  'sd62045;
    data[3014] = -'sd17457;
    data[3015] =  'sd76556;
    data[3016] =  'sd55098;
    data[3017] = -'sd52192;
    data[3018] =  'sd66722;
    data[3019] =  'sd5928;
    data[3020] =  'sd29640;
    data[3021] = -'sd15641;
    data[3022] = -'sd78205;
    data[3023] = -'sd63343;
    data[3024] =  'sd10967;
    data[3025] =  'sd54835;
    data[3026] = -'sd53507;
    data[3027] =  'sd60147;
    data[3028] = -'sd26947;
    data[3029] =  'sd29106;
    data[3030] = -'sd18311;
    data[3031] =  'sd72286;
    data[3032] =  'sd33748;
    data[3033] =  'sd4899;
    data[3034] =  'sd24495;
    data[3035] = -'sd41366;
    data[3036] = -'sd42989;
    data[3037] = -'sd51104;
    data[3038] =  'sd72162;
    data[3039] =  'sd33128;
    data[3040] =  'sd1799;
    data[3041] =  'sd8995;
    data[3042] =  'sd44975;
    data[3043] =  'sd61034;
    data[3044] = -'sd22512;
    data[3045] =  'sd51281;
    data[3046] = -'sd71277;
    data[3047] = -'sd28703;
    data[3048] =  'sd20326;
    data[3049] = -'sd62211;
    data[3050] =  'sd16627;
    data[3051] = -'sd80706;
    data[3052] = -'sd75848;
    data[3053] = -'sd51558;
    data[3054] =  'sd69892;
    data[3055] =  'sd21778;
    data[3056] = -'sd54951;
    data[3057] =  'sd52927;
    data[3058] = -'sd63047;
    data[3059] =  'sd12447;
    data[3060] =  'sd62235;
    data[3061] = -'sd16507;
    data[3062] =  'sd81306;
    data[3063] =  'sd78848;
    data[3064] =  'sd66558;
    data[3065] =  'sd5108;
    data[3066] =  'sd25540;
    data[3067] = -'sd36141;
    data[3068] = -'sd16864;
    data[3069] =  'sd79521;
    data[3070] =  'sd69923;
    data[3071] =  'sd21933;
    data[3072] = -'sd54176;
    data[3073] =  'sd56802;
    data[3074] = -'sd43672;
    data[3075] = -'sd54519;
    data[3076] =  'sd55087;
    data[3077] = -'sd52247;
    data[3078] =  'sd66447;
    data[3079] =  'sd4553;
    data[3080] =  'sd22765;
    data[3081] = -'sd50016;
    data[3082] =  'sd77602;
    data[3083] =  'sd60328;
    data[3084] = -'sd26042;
    data[3085] =  'sd33631;
    data[3086] =  'sd4314;
    data[3087] =  'sd21570;
    data[3088] = -'sd55991;
    data[3089] =  'sd47727;
    data[3090] =  'sd74794;
    data[3091] =  'sd46288;
    data[3092] =  'sd67599;
    data[3093] =  'sd10313;
    data[3094] =  'sd51565;
    data[3095] = -'sd69857;
    data[3096] = -'sd21603;
    data[3097] =  'sd55826;
    data[3098] = -'sd48552;
    data[3099] = -'sd78919;
    data[3100] = -'sd66913;
    data[3101] = -'sd6883;
    data[3102] = -'sd34415;
    data[3103] = -'sd8234;
    data[3104] = -'sd41170;
    data[3105] = -'sd42009;
    data[3106] = -'sd46204;
    data[3107] = -'sd67179;
    data[3108] = -'sd8213;
    data[3109] = -'sd41065;
    data[3110] = -'sd41484;
    data[3111] = -'sd43579;
    data[3112] = -'sd54054;
    data[3113] =  'sd57412;
    data[3114] = -'sd40622;
    data[3115] = -'sd39269;
    data[3116] = -'sd32504;
    data[3117] =  'sd1321;
    data[3118] =  'sd6605;
    data[3119] =  'sd33025;
    data[3120] =  'sd1284;
    data[3121] =  'sd6420;
    data[3122] =  'sd32100;
    data[3123] = -'sd3341;
    data[3124] = -'sd16705;
    data[3125] =  'sd80316;
    data[3126] =  'sd73898;
    data[3127] =  'sd41808;
    data[3128] =  'sd45199;
    data[3129] =  'sd62154;
    data[3130] = -'sd16912;
    data[3131] =  'sd79281;
    data[3132] =  'sd68723;
    data[3133] =  'sd15933;
    data[3134] =  'sd79665;
    data[3135] =  'sd70643;
    data[3136] =  'sd25533;
    data[3137] = -'sd36176;
    data[3138] = -'sd17039;
    data[3139] =  'sd78646;
    data[3140] =  'sd65548;
    data[3141] =  'sd58;
    data[3142] =  'sd290;
    data[3143] =  'sd1450;
    data[3144] =  'sd7250;
    data[3145] =  'sd36250;
    data[3146] =  'sd17409;
    data[3147] = -'sd76796;
    data[3148] = -'sd56298;
    data[3149] =  'sd46192;
    data[3150] =  'sd67119;
    data[3151] =  'sd7913;
    data[3152] =  'sd39565;
    data[3153] =  'sd33984;
    data[3154] =  'sd6079;
    data[3155] =  'sd30395;
    data[3156] = -'sd11866;
    data[3157] = -'sd59330;
    data[3158] =  'sd31032;
    data[3159] = -'sd8681;
    data[3160] = -'sd43405;
    data[3161] = -'sd53184;
    data[3162] =  'sd61762;
    data[3163] = -'sd18872;
    data[3164] =  'sd69481;
    data[3165] =  'sd19723;
    data[3166] = -'sd65226;
    data[3167] =  'sd1552;
    data[3168] =  'sd7760;
    data[3169] =  'sd38800;
    data[3170] =  'sd30159;
    data[3171] = -'sd13046;
    data[3172] = -'sd65230;
    data[3173] =  'sd1532;
    data[3174] =  'sd7660;
    data[3175] =  'sd38300;
    data[3176] =  'sd27659;
    data[3177] = -'sd25546;
    data[3178] =  'sd36111;
    data[3179] =  'sd16714;
    data[3180] = -'sd80271;
    data[3181] = -'sd73673;
    data[3182] = -'sd40683;
    data[3183] = -'sd39574;
    data[3184] = -'sd34029;
    data[3185] = -'sd6304;
    data[3186] = -'sd31520;
    data[3187] =  'sd6241;
    data[3188] =  'sd31205;
    data[3189] = -'sd7816;
    data[3190] = -'sd39080;
    data[3191] = -'sd31559;
    data[3192] =  'sd6046;
    data[3193] =  'sd30230;
    data[3194] = -'sd12691;
    data[3195] = -'sd63455;
    data[3196] =  'sd10407;
    data[3197] =  'sd52035;
    data[3198] = -'sd67507;
    data[3199] = -'sd9853;
    data[3200] = -'sd49265;
    data[3201] =  'sd81357;
    data[3202] =  'sd79103;
    data[3203] =  'sd67833;
    data[3204] =  'sd11483;
    data[3205] =  'sd57415;
    data[3206] = -'sd40607;
    data[3207] = -'sd39194;
    data[3208] = -'sd32129;
    data[3209] =  'sd3196;
    data[3210] =  'sd15980;
    data[3211] =  'sd79900;
    data[3212] =  'sd71818;
    data[3213] =  'sd31408;
    data[3214] = -'sd6801;
    data[3215] = -'sd34005;
    data[3216] = -'sd6184;
    data[3217] = -'sd30920;
    data[3218] =  'sd9241;
    data[3219] =  'sd46205;
    data[3220] =  'sd67184;
    data[3221] =  'sd8238;
    data[3222] =  'sd41190;
    data[3223] =  'sd42109;
    data[3224] =  'sd46704;
    data[3225] =  'sd69679;
    data[3226] =  'sd20713;
    data[3227] = -'sd60276;
    data[3228] =  'sd26302;
    data[3229] = -'sd32331;
    data[3230] =  'sd2186;
    data[3231] =  'sd10930;
    data[3232] =  'sd54650;
    data[3233] = -'sd54432;
    data[3234] =  'sd55522;
    data[3235] = -'sd50072;
    data[3236] =  'sd77322;
    data[3237] =  'sd58928;
    data[3238] = -'sd33042;
    data[3239] = -'sd1369;
    data[3240] = -'sd6845;
    data[3241] = -'sd34225;
    data[3242] = -'sd7284;
    data[3243] = -'sd36420;
    data[3244] = -'sd18259;
    data[3245] =  'sd72546;
    data[3246] =  'sd35048;
    data[3247] =  'sd11399;
    data[3248] =  'sd56995;
    data[3249] = -'sd42707;
    data[3250] = -'sd49694;
    data[3251] =  'sd79212;
    data[3252] =  'sd68378;
    data[3253] =  'sd14208;
    data[3254] =  'sd71040;
    data[3255] =  'sd27518;
    data[3256] = -'sd26251;
    data[3257] =  'sd32586;
    data[3258] = -'sd911;
    data[3259] = -'sd4555;
    data[3260] = -'sd22775;
    data[3261] =  'sd49966;
    data[3262] = -'sd77852;
    data[3263] = -'sd61578;
    data[3264] =  'sd19792;
    data[3265] = -'sd64881;
    data[3266] =  'sd3277;
    data[3267] =  'sd16385;
    data[3268] = -'sd81916;
    data[3269] = -'sd81898;
    data[3270] = -'sd81808;
    data[3271] = -'sd81358;
    data[3272] = -'sd79108;
    data[3273] = -'sd67858;
    data[3274] = -'sd11608;
    data[3275] = -'sd58040;
    data[3276] =  'sd37482;
    data[3277] =  'sd23569;
    data[3278] = -'sd45996;
    data[3279] = -'sd66139;
    data[3280] = -'sd3013;
    data[3281] = -'sd15065;
    data[3282] = -'sd75325;
    data[3283] = -'sd48943;
    data[3284] = -'sd80874;
    data[3285] = -'sd76688;
    data[3286] = -'sd55758;
    data[3287] =  'sd48892;
    data[3288] =  'sd80619;
    data[3289] =  'sd75413;
    data[3290] =  'sd49383;
    data[3291] = -'sd80767;
    data[3292] = -'sd76153;
    data[3293] = -'sd53083;
    data[3294] =  'sd62267;
    data[3295] = -'sd16347;
    data[3296] = -'sd81735;
    data[3297] = -'sd80993;
    data[3298] = -'sd77283;
    data[3299] = -'sd58733;
    data[3300] =  'sd34017;
    data[3301] =  'sd6244;
    data[3302] =  'sd31220;
    data[3303] = -'sd7741;
    data[3304] = -'sd38705;
    data[3305] = -'sd29684;
    data[3306] =  'sd15421;
    data[3307] =  'sd77105;
    data[3308] =  'sd57843;
    data[3309] = -'sd38467;
    data[3310] = -'sd28494;
    data[3311] =  'sd21371;
    data[3312] = -'sd56986;
    data[3313] =  'sd42752;
    data[3314] =  'sd49919;
    data[3315] = -'sd78087;
    data[3316] = -'sd62753;
    data[3317] =  'sd13917;
    data[3318] =  'sd69585;
    data[3319] =  'sd20243;
    data[3320] = -'sd62626;
    data[3321] =  'sd14552;
    data[3322] =  'sd72760;
    data[3323] =  'sd36118;
    data[3324] =  'sd16749;
    data[3325] = -'sd80096;
    data[3326] = -'sd72798;
    data[3327] = -'sd36308;
    data[3328] = -'sd17699;
    data[3329] =  'sd75346;
    data[3330] =  'sd49048;
    data[3331] =  'sd81399;
    data[3332] =  'sd79313;
    data[3333] =  'sd68883;
    data[3334] =  'sd16733;
    data[3335] = -'sd80176;
    data[3336] = -'sd73198;
    data[3337] = -'sd38308;
    data[3338] = -'sd27699;
    data[3339] =  'sd25346;
    data[3340] = -'sd37111;
    data[3341] = -'sd21714;
    data[3342] =  'sd55271;
    data[3343] = -'sd51327;
    data[3344] =  'sd71047;
    data[3345] =  'sd27553;
    data[3346] = -'sd26076;
    data[3347] =  'sd33461;
    data[3348] =  'sd3464;
    data[3349] =  'sd17320;
    data[3350] = -'sd77241;
    data[3351] = -'sd58523;
    data[3352] =  'sd35067;
    data[3353] =  'sd11494;
    data[3354] =  'sd57470;
    data[3355] = -'sd40332;
    data[3356] = -'sd37819;
    data[3357] = -'sd25254;
    data[3358] =  'sd37571;
    data[3359] =  'sd24014;
    data[3360] = -'sd43771;
    data[3361] = -'sd55014;
    data[3362] =  'sd52612;
    data[3363] = -'sd64622;
    data[3364] =  'sd4572;
    data[3365] =  'sd22860;
    data[3366] = -'sd49541;
    data[3367] =  'sd79977;
    data[3368] =  'sd72203;
    data[3369] =  'sd33333;
    data[3370] =  'sd2824;
    data[3371] =  'sd14120;
    data[3372] =  'sd70600;
    data[3373] =  'sd25318;
    data[3374] = -'sd37251;
    data[3375] = -'sd22414;
    data[3376] =  'sd51771;
    data[3377] = -'sd68827;
    data[3378] = -'sd16453;
    data[3379] =  'sd81576;
    data[3380] =  'sd80198;
    data[3381] =  'sd73308;
    data[3382] =  'sd38858;
    data[3383] =  'sd30449;
    data[3384] = -'sd11596;
    data[3385] = -'sd57980;
    data[3386] =  'sd37782;
    data[3387] =  'sd25069;
    data[3388] = -'sd38496;
    data[3389] = -'sd28639;
    data[3390] =  'sd20646;
    data[3391] = -'sd60611;
    data[3392] =  'sd24627;
    data[3393] = -'sd40706;
    data[3394] = -'sd39689;
    data[3395] = -'sd34604;
    data[3396] = -'sd9179;
    data[3397] = -'sd45895;
    data[3398] = -'sd65634;
    data[3399] = -'sd488;
    data[3400] = -'sd2440;
    data[3401] = -'sd12200;
    data[3402] = -'sd61000;
    data[3403] =  'sd22682;
    data[3404] = -'sd50431;
    data[3405] =  'sd75527;
    data[3406] =  'sd49953;
    data[3407] = -'sd77917;
    data[3408] = -'sd61903;
    data[3409] =  'sd18167;
    data[3410] = -'sd73006;
    data[3411] = -'sd37348;
    data[3412] = -'sd22899;
    data[3413] =  'sd49346;
    data[3414] = -'sd80952;
    data[3415] = -'sd77078;
    data[3416] = -'sd57708;
    data[3417] =  'sd39142;
    data[3418] =  'sd31869;
    data[3419] = -'sd4496;
    data[3420] = -'sd22480;
    data[3421] =  'sd51441;
    data[3422] = -'sd70477;
    data[3423] = -'sd24703;
    data[3424] =  'sd40326;
    data[3425] =  'sd37789;
    data[3426] =  'sd25104;
    data[3427] = -'sd38321;
    data[3428] = -'sd27764;
    data[3429] =  'sd25021;
    data[3430] = -'sd38736;
    data[3431] = -'sd29839;
    data[3432] =  'sd14646;
    data[3433] =  'sd73230;
    data[3434] =  'sd38468;
    data[3435] =  'sd28499;
    data[3436] = -'sd21346;
    data[3437] =  'sd57111;
    data[3438] = -'sd42127;
    data[3439] = -'sd46794;
    data[3440] = -'sd70129;
    data[3441] = -'sd22963;
    data[3442] =  'sd49026;
    data[3443] =  'sd81289;
    data[3444] =  'sd78763;
    data[3445] =  'sd66133;
    data[3446] =  'sd2983;
    data[3447] =  'sd14915;
    data[3448] =  'sd74575;
    data[3449] =  'sd45193;
    data[3450] =  'sd62124;
    data[3451] = -'sd17062;
    data[3452] =  'sd78531;
    data[3453] =  'sd64973;
    data[3454] = -'sd2817;
    data[3455] = -'sd14085;
    data[3456] = -'sd70425;
    data[3457] = -'sd24443;
    data[3458] =  'sd41626;
    data[3459] =  'sd44289;
    data[3460] =  'sd57604;
    data[3461] = -'sd39662;
    data[3462] = -'sd34469;
    data[3463] = -'sd8504;
    data[3464] = -'sd42520;
    data[3465] = -'sd48759;
    data[3466] = -'sd79954;
    data[3467] = -'sd72088;
    data[3468] = -'sd32758;
    data[3469] =  'sd51;
    data[3470] =  'sd255;
    data[3471] =  'sd1275;
    data[3472] =  'sd6375;
    data[3473] =  'sd31875;
    data[3474] = -'sd4466;
    data[3475] = -'sd22330;
    data[3476] =  'sd52191;
    data[3477] = -'sd66727;
    data[3478] = -'sd5953;
    data[3479] = -'sd29765;
    data[3480] =  'sd15016;
    data[3481] =  'sd75080;
    data[3482] =  'sd47718;
    data[3483] =  'sd74749;
    data[3484] =  'sd46063;
    data[3485] =  'sd66474;
    data[3486] =  'sd4688;
    data[3487] =  'sd23440;
    data[3488] = -'sd46641;
    data[3489] = -'sd69364;
    data[3490] = -'sd19138;
    data[3491] =  'sd68151;
    data[3492] =  'sd13073;
    data[3493] =  'sd65365;
    data[3494] = -'sd857;
    data[3495] = -'sd4285;
    data[3496] = -'sd21425;
    data[3497] =  'sd56716;
    data[3498] = -'sd44102;
    data[3499] = -'sd56669;
    data[3500] =  'sd44337;
    data[3501] =  'sd57844;
    data[3502] = -'sd38462;
    data[3503] = -'sd28469;
    data[3504] =  'sd21496;
    data[3505] = -'sd56361;
    data[3506] =  'sd45877;
    data[3507] =  'sd65544;
    data[3508] =  'sd38;
    data[3509] =  'sd190;
    data[3510] =  'sd950;
    data[3511] =  'sd4750;
    data[3512] =  'sd23750;
    data[3513] = -'sd45091;
    data[3514] = -'sd61614;
    data[3515] =  'sd19612;
    data[3516] = -'sd65781;
    data[3517] = -'sd1223;
    data[3518] = -'sd6115;
    data[3519] = -'sd30575;
    data[3520] =  'sd10966;
    data[3521] =  'sd54830;
    data[3522] = -'sd53532;
    data[3523] =  'sd60022;
    data[3524] = -'sd27572;
    data[3525] =  'sd25981;
    data[3526] = -'sd33936;
    data[3527] = -'sd5839;
    data[3528] = -'sd29195;
    data[3529] =  'sd17866;
    data[3530] = -'sd74511;
    data[3531] = -'sd44873;
    data[3532] = -'sd60524;
    data[3533] =  'sd25062;
    data[3534] = -'sd38531;
    data[3535] = -'sd28814;
    data[3536] =  'sd19771;
    data[3537] = -'sd64986;
    data[3538] =  'sd2752;
    data[3539] =  'sd13760;
    data[3540] =  'sd68800;
    data[3541] =  'sd16318;
    data[3542] =  'sd81590;
    data[3543] =  'sd80268;
    data[3544] =  'sd73658;
    data[3545] =  'sd40608;
    data[3546] =  'sd39199;
    data[3547] =  'sd32154;
    data[3548] = -'sd3071;
    data[3549] = -'sd15355;
    data[3550] = -'sd76775;
    data[3551] = -'sd56193;
    data[3552] =  'sd46717;
    data[3553] =  'sd69744;
    data[3554] =  'sd21038;
    data[3555] = -'sd58651;
    data[3556] =  'sd34427;
    data[3557] =  'sd8294;
    data[3558] =  'sd41470;
    data[3559] =  'sd43509;
    data[3560] =  'sd53704;
    data[3561] = -'sd59162;
    data[3562] =  'sd31872;
    data[3563] = -'sd4481;
    data[3564] = -'sd22405;
    data[3565] =  'sd51816;
    data[3566] = -'sd68602;
    data[3567] = -'sd15328;
    data[3568] = -'sd76640;
    data[3569] = -'sd55518;
    data[3570] =  'sd50092;
    data[3571] = -'sd77222;
    data[3572] = -'sd58428;
    data[3573] =  'sd35542;
    data[3574] =  'sd13869;
    data[3575] =  'sd69345;
    data[3576] =  'sd19043;
    data[3577] = -'sd68626;
    data[3578] = -'sd15448;
    data[3579] = -'sd77240;
    data[3580] = -'sd58518;
    data[3581] =  'sd35092;
    data[3582] =  'sd11619;
    data[3583] =  'sd58095;
    data[3584] = -'sd37207;
    data[3585] = -'sd22194;
    data[3586] =  'sd52871;
    data[3587] = -'sd63327;
    data[3588] =  'sd11047;
    data[3589] =  'sd55235;
    data[3590] = -'sd51507;
    data[3591] =  'sd70147;
    data[3592] =  'sd23053;
    data[3593] = -'sd48576;
    data[3594] = -'sd79039;
    data[3595] = -'sd67513;
    data[3596] = -'sd9883;
    data[3597] = -'sd49415;
    data[3598] =  'sd80607;
    data[3599] =  'sd75353;
    data[3600] =  'sd49083;
    data[3601] =  'sd81574;
    data[3602] =  'sd80188;
    data[3603] =  'sd73258;
    data[3604] =  'sd38608;
    data[3605] =  'sd29199;
    data[3606] = -'sd17846;
    data[3607] =  'sd74611;
    data[3608] =  'sd45373;
    data[3609] =  'sd63024;
    data[3610] = -'sd12562;
    data[3611] = -'sd62810;
    data[3612] =  'sd13632;
    data[3613] =  'sd68160;
    data[3614] =  'sd13118;
    data[3615] =  'sd65590;
    data[3616] =  'sd268;
    data[3617] =  'sd1340;
    data[3618] =  'sd6700;
    data[3619] =  'sd33500;
    data[3620] =  'sd3659;
    data[3621] =  'sd18295;
    data[3622] = -'sd72366;
    data[3623] = -'sd34148;
    data[3624] = -'sd6899;
    data[3625] = -'sd34495;
    data[3626] = -'sd8634;
    data[3627] = -'sd43170;
    data[3628] = -'sd52009;
    data[3629] =  'sd67637;
    data[3630] =  'sd10503;
    data[3631] =  'sd52515;
    data[3632] = -'sd65107;
    data[3633] =  'sd2147;
    data[3634] =  'sd10735;
    data[3635] =  'sd53675;
    data[3636] = -'sd59307;
    data[3637] =  'sd31147;
    data[3638] = -'sd8106;
    data[3639] = -'sd40530;
    data[3640] = -'sd38809;
    data[3641] = -'sd30204;
    data[3642] =  'sd12821;
    data[3643] =  'sd64105;
    data[3644] = -'sd7157;
    data[3645] = -'sd35785;
    data[3646] = -'sd15084;
    data[3647] = -'sd75420;
    data[3648] = -'sd49418;
    data[3649] =  'sd80592;
    data[3650] =  'sd75278;
    data[3651] =  'sd48708;
    data[3652] =  'sd79699;
    data[3653] =  'sd70813;
    data[3654] =  'sd26383;
    data[3655] = -'sd31926;
    data[3656] =  'sd4211;
    data[3657] =  'sd21055;
    data[3658] = -'sd58566;
    data[3659] =  'sd34852;
    data[3660] =  'sd10419;
    data[3661] =  'sd52095;
    data[3662] = -'sd67207;
    data[3663] = -'sd8353;
    data[3664] = -'sd41765;
    data[3665] = -'sd44984;
    data[3666] = -'sd61079;
    data[3667] =  'sd22287;
    data[3668] = -'sd52406;
    data[3669] =  'sd65652;
    data[3670] =  'sd578;
    data[3671] =  'sd2890;
    data[3672] =  'sd14450;
    data[3673] =  'sd72250;
    data[3674] =  'sd33568;
    data[3675] =  'sd3999;
    data[3676] =  'sd19995;
    data[3677] = -'sd63866;
    data[3678] =  'sd8352;
    data[3679] =  'sd41760;
    data[3680] =  'sd44959;
    data[3681] =  'sd60954;
    data[3682] = -'sd22912;
    data[3683] =  'sd49281;
    data[3684] = -'sd81277;
    data[3685] = -'sd78703;
    data[3686] = -'sd65833;
    data[3687] = -'sd1483;
    data[3688] = -'sd7415;
    data[3689] = -'sd37075;
    data[3690] = -'sd21534;
    data[3691] =  'sd56171;
    data[3692] = -'sd46827;
    data[3693] = -'sd70294;
    data[3694] = -'sd23788;
    data[3695] =  'sd44901;
    data[3696] =  'sd60664;
    data[3697] = -'sd24362;
    data[3698] =  'sd42031;
    data[3699] =  'sd46314;
    data[3700] =  'sd67729;
    data[3701] =  'sd10963;
    data[3702] =  'sd54815;
    data[3703] = -'sd53607;
    data[3704] =  'sd59647;
    data[3705] = -'sd29447;
    data[3706] =  'sd16606;
    data[3707] = -'sd80811;
    data[3708] = -'sd76373;
    data[3709] = -'sd54183;
    data[3710] =  'sd56767;
    data[3711] = -'sd43847;
    data[3712] = -'sd55394;
    data[3713] =  'sd50712;
    data[3714] = -'sd74122;
    data[3715] = -'sd42928;
    data[3716] = -'sd50799;
    data[3717] =  'sd73687;
    data[3718] =  'sd40753;
    data[3719] =  'sd39924;
    data[3720] =  'sd35779;
    data[3721] =  'sd15054;
    data[3722] =  'sd75270;
    data[3723] =  'sd48668;
    data[3724] =  'sd79499;
    data[3725] =  'sd69813;
    data[3726] =  'sd21383;
    data[3727] = -'sd56926;
    data[3728] =  'sd43052;
    data[3729] =  'sd51419;
    data[3730] = -'sd70587;
    data[3731] = -'sd25253;
    data[3732] =  'sd37576;
    data[3733] =  'sd24039;
    data[3734] = -'sd43646;
    data[3735] = -'sd54389;
    data[3736] =  'sd55737;
    data[3737] = -'sd48997;
    data[3738] = -'sd81144;
    data[3739] = -'sd78038;
    data[3740] = -'sd62508;
    data[3741] =  'sd15142;
    data[3742] =  'sd75710;
    data[3743] =  'sd50868;
    data[3744] = -'sd73342;
    data[3745] = -'sd39028;
    data[3746] = -'sd31299;
    data[3747] =  'sd7346;
    data[3748] =  'sd36730;
    data[3749] =  'sd19809;
    data[3750] = -'sd64796;
    data[3751] =  'sd3702;
    data[3752] =  'sd18510;
    data[3753] = -'sd71291;
    data[3754] = -'sd28773;
    data[3755] =  'sd19976;
    data[3756] = -'sd63961;
    data[3757] =  'sd7877;
    data[3758] =  'sd39385;
    data[3759] =  'sd33084;
    data[3760] =  'sd1579;
    data[3761] =  'sd7895;
    data[3762] =  'sd39475;
    data[3763] =  'sd33534;
    data[3764] =  'sd3829;
    data[3765] =  'sd19145;
    data[3766] = -'sd68116;
    data[3767] = -'sd12898;
    data[3768] = -'sd64490;
    data[3769] =  'sd5232;
    data[3770] =  'sd26160;
    data[3771] = -'sd33041;
    data[3772] = -'sd1364;
    data[3773] = -'sd6820;
    data[3774] = -'sd34100;
    data[3775] = -'sd6659;
    data[3776] = -'sd33295;
    data[3777] = -'sd2634;
    data[3778] = -'sd13170;
    data[3779] = -'sd65850;
    data[3780] = -'sd1568;
    data[3781] = -'sd7840;
    data[3782] = -'sd39200;
    data[3783] = -'sd32159;
    data[3784] =  'sd3046;
    data[3785] =  'sd15230;
    data[3786] =  'sd76150;
    data[3787] =  'sd53068;
    data[3788] = -'sd62342;
    data[3789] =  'sd15972;
    data[3790] =  'sd79860;
    data[3791] =  'sd71618;
    data[3792] =  'sd30408;
    data[3793] = -'sd11801;
    data[3794] = -'sd59005;
    data[3795] =  'sd32657;
    data[3796] = -'sd556;
    data[3797] = -'sd2780;
    data[3798] = -'sd13900;
    data[3799] = -'sd69500;
    data[3800] = -'sd19818;
    data[3801] =  'sd64751;
    data[3802] = -'sd3927;
    data[3803] = -'sd19635;
    data[3804] =  'sd65666;
    data[3805] =  'sd648;
    data[3806] =  'sd3240;
    data[3807] =  'sd16200;
    data[3808] =  'sd81000;
    data[3809] =  'sd77318;
    data[3810] =  'sd58908;
    data[3811] = -'sd33142;
    data[3812] = -'sd1869;
    data[3813] = -'sd9345;
    data[3814] = -'sd46725;
    data[3815] = -'sd69784;
    data[3816] = -'sd21238;
    data[3817] =  'sd57651;
    data[3818] = -'sd39427;
    data[3819] = -'sd33294;
    data[3820] = -'sd2629;
    data[3821] = -'sd13145;
    data[3822] = -'sd65725;
    data[3823] = -'sd943;
    data[3824] = -'sd4715;
    data[3825] = -'sd23575;
    data[3826] =  'sd45966;
    data[3827] =  'sd65989;
    data[3828] =  'sd2263;
    data[3829] =  'sd11315;
    data[3830] =  'sd56575;
    data[3831] = -'sd44807;
    data[3832] = -'sd60194;
    data[3833] =  'sd26712;
    data[3834] = -'sd30281;
    data[3835] =  'sd12436;
    data[3836] =  'sd62180;
    data[3837] = -'sd16782;
    data[3838] =  'sd79931;
    data[3839] =  'sd71973;
    data[3840] =  'sd32183;
    data[3841] = -'sd2926;
    data[3842] = -'sd14630;
    data[3843] = -'sd73150;
    data[3844] = -'sd38068;
    data[3845] = -'sd26499;
    data[3846] =  'sd31346;
    data[3847] = -'sd7111;
    data[3848] = -'sd35555;
    data[3849] = -'sd13934;
    data[3850] = -'sd69670;
    data[3851] = -'sd20668;
    data[3852] =  'sd60501;
    data[3853] = -'sd25177;
    data[3854] =  'sd37956;
    data[3855] =  'sd25939;
    data[3856] = -'sd34146;
    data[3857] = -'sd6889;
    data[3858] = -'sd34445;
    data[3859] = -'sd8384;
    data[3860] = -'sd41920;
    data[3861] = -'sd45759;
    data[3862] = -'sd64954;
    data[3863] =  'sd2912;
    data[3864] =  'sd14560;
    data[3865] =  'sd72800;
    data[3866] =  'sd36318;
    data[3867] =  'sd17749;
    data[3868] = -'sd75096;
    data[3869] = -'sd47798;
    data[3870] = -'sd75149;
    data[3871] = -'sd48063;
    data[3872] = -'sd76474;
    data[3873] = -'sd54688;
    data[3874] =  'sd54242;
    data[3875] = -'sd56472;
    data[3876] =  'sd45322;
    data[3877] =  'sd62769;
    data[3878] = -'sd13837;
    data[3879] = -'sd69185;
    data[3880] = -'sd18243;
    data[3881] =  'sd72626;
    data[3882] =  'sd35448;
    data[3883] =  'sd13399;
    data[3884] =  'sd66995;
    data[3885] =  'sd7293;
    data[3886] =  'sd36465;
    data[3887] =  'sd18484;
    data[3888] = -'sd71421;
    data[3889] = -'sd29423;
    data[3890] =  'sd16726;
    data[3891] = -'sd80211;
    data[3892] = -'sd73373;
    data[3893] = -'sd39183;
    data[3894] = -'sd32074;
    data[3895] =  'sd3471;
    data[3896] =  'sd17355;
    data[3897] = -'sd77066;
    data[3898] = -'sd57648;
    data[3899] =  'sd39442;
    data[3900] =  'sd33369;
    data[3901] =  'sd3004;
    data[3902] =  'sd15020;
    data[3903] =  'sd75100;
    data[3904] =  'sd47818;
    data[3905] =  'sd75249;
    data[3906] =  'sd48563;
    data[3907] =  'sd78974;
    data[3908] =  'sd67188;
    data[3909] =  'sd8258;
    data[3910] =  'sd41290;
    data[3911] =  'sd42609;
    data[3912] =  'sd49204;
    data[3913] = -'sd81662;
    data[3914] = -'sd80628;
    data[3915] = -'sd75458;
    data[3916] = -'sd49608;
    data[3917] =  'sd79642;
    data[3918] =  'sd70528;
    data[3919] =  'sd24958;
    data[3920] = -'sd39051;
    data[3921] = -'sd31414;
    data[3922] =  'sd6771;
    data[3923] =  'sd33855;
    data[3924] =  'sd5434;
    data[3925] =  'sd27170;
    data[3926] = -'sd27991;
    data[3927] =  'sd23886;
    data[3928] = -'sd44411;
    data[3929] = -'sd58214;
    data[3930] =  'sd36612;
    data[3931] =  'sd19219;
    data[3932] = -'sd67746;
    data[3933] = -'sd11048;
    data[3934] = -'sd55240;
    data[3935] =  'sd51482;
    data[3936] = -'sd70272;
    data[3937] = -'sd23678;
    data[3938] =  'sd45451;
    data[3939] =  'sd63414;
    data[3940] = -'sd10612;
    data[3941] = -'sd53060;
    data[3942] =  'sd62382;
    data[3943] = -'sd15772;
    data[3944] = -'sd78860;
    data[3945] = -'sd66618;
    data[3946] = -'sd5408;
    data[3947] = -'sd27040;
    data[3948] =  'sd28641;
    data[3949] = -'sd20636;
    data[3950] =  'sd60661;
    data[3951] = -'sd24377;
    data[3952] =  'sd41956;
    data[3953] =  'sd45939;
    data[3954] =  'sd65854;
    data[3955] =  'sd1588;
    data[3956] =  'sd7940;
    data[3957] =  'sd39700;
    data[3958] =  'sd34659;
    data[3959] =  'sd9454;
    data[3960] =  'sd47270;
    data[3961] =  'sd72509;
    data[3962] =  'sd34863;
    data[3963] =  'sd10474;
    data[3964] =  'sd52370;
    data[3965] = -'sd65832;
    data[3966] = -'sd1478;
    data[3967] = -'sd7390;
    data[3968] = -'sd36950;
    data[3969] = -'sd20909;
    data[3970] =  'sd59296;
    data[3971] = -'sd31202;
    data[3972] =  'sd7831;
    data[3973] =  'sd39155;
    data[3974] =  'sd31934;
    data[3975] = -'sd4171;
    data[3976] = -'sd20855;
    data[3977] =  'sd59566;
    data[3978] = -'sd29852;
    data[3979] =  'sd14581;
    data[3980] =  'sd72905;
    data[3981] =  'sd36843;
    data[3982] =  'sd20374;
    data[3983] = -'sd61971;
    data[3984] =  'sd17827;
    data[3985] = -'sd74706;
    data[3986] = -'sd45848;
    data[3987] = -'sd65399;
    data[3988] =  'sd687;
    data[3989] =  'sd3435;
    data[3990] =  'sd17175;
    data[3991] = -'sd77966;
    data[3992] = -'sd62148;
    data[3993] =  'sd16942;
    data[3994] = -'sd79131;
    data[3995] = -'sd67973;
    data[3996] = -'sd12183;
    data[3997] = -'sd60915;
    data[3998] =  'sd23107;
    data[3999] = -'sd48306;
    data[4000] = -'sd77689;
    data[4001] = -'sd60763;
    data[4002] =  'sd23867;
    data[4003] = -'sd44506;
    data[4004] = -'sd58689;
    data[4005] =  'sd34237;
    data[4006] =  'sd7344;
    data[4007] =  'sd36720;
    data[4008] =  'sd19759;
    data[4009] = -'sd65046;
    data[4010] =  'sd2452;
    data[4011] =  'sd12260;
    data[4012] =  'sd61300;
    data[4013] = -'sd21182;
    data[4014] =  'sd57931;
    data[4015] = -'sd38027;
    data[4016] = -'sd26294;
    data[4017] =  'sd32371;
    data[4018] = -'sd1986;
    data[4019] = -'sd9930;
    data[4020] = -'sd49650;
    data[4021] =  'sd79432;
    data[4022] =  'sd69478;
    data[4023] =  'sd19708;
    data[4024] = -'sd65301;
    data[4025] =  'sd1177;
    data[4026] =  'sd5885;
    data[4027] =  'sd29425;
    data[4028] = -'sd16716;
    data[4029] =  'sd80261;
    data[4030] =  'sd73623;
    data[4031] =  'sd40433;
    data[4032] =  'sd38324;
    data[4033] =  'sd27779;
    data[4034] = -'sd24946;
    data[4035] =  'sd39111;
    data[4036] =  'sd31714;
    data[4037] = -'sd5271;
    data[4038] = -'sd26355;
    data[4039] =  'sd32066;
    data[4040] = -'sd3511;
    data[4041] = -'sd17555;
    data[4042] =  'sd76066;
    data[4043] =  'sd52648;
    data[4044] = -'sd64442;
    data[4045] =  'sd5472;
    data[4046] =  'sd27360;
    data[4047] = -'sd27041;
    data[4048] =  'sd28636;
    data[4049] = -'sd20661;
    data[4050] =  'sd60536;
    data[4051] = -'sd25002;
    data[4052] =  'sd38831;
    data[4053] =  'sd30314;
    data[4054] = -'sd12271;
    data[4055] = -'sd61355;
    data[4056] =  'sd20907;
    data[4057] = -'sd59306;
    data[4058] =  'sd31152;
    data[4059] = -'sd8081;
    data[4060] = -'sd40405;
    data[4061] = -'sd38184;
    data[4062] = -'sd27079;
    data[4063] =  'sd28446;
    data[4064] = -'sd21611;
    data[4065] =  'sd55786;
    data[4066] = -'sd48752;
    data[4067] = -'sd79919;
    data[4068] = -'sd71913;
    data[4069] = -'sd31883;
    data[4070] =  'sd4426;
    data[4071] =  'sd22130;
    data[4072] = -'sd53191;
    data[4073] =  'sd61727;
    data[4074] = -'sd19047;
    data[4075] =  'sd68606;
    data[4076] =  'sd15348;
    data[4077] =  'sd76740;
    data[4078] =  'sd56018;
    data[4079] = -'sd47592;
    data[4080] = -'sd74119;
    data[4081] = -'sd42913;
    data[4082] = -'sd50724;
    data[4083] =  'sd74062;
    data[4084] =  'sd42628;
    data[4085] =  'sd49299;
    data[4086] = -'sd81187;
    data[4087] = -'sd78253;
    data[4088] = -'sd63583;
    data[4089] =  'sd9767;
    data[4090] =  'sd48835;
    data[4091] =  'sd80334;
    data[4092] =  'sd73988;
    data[4093] =  'sd42258;
    data[4094] =  'sd47449;
    data[4095] =  'sd73404;
    data[4096] =  'sd39338;
    data[4097] =  'sd32849;
    data[4098] =  'sd404;
    data[4099] =  'sd2020;
    data[4100] =  'sd10100;
    data[4101] =  'sd50500;
    data[4102] = -'sd75182;
    data[4103] = -'sd48228;
    data[4104] = -'sd77299;
    data[4105] = -'sd58813;
    data[4106] =  'sd33617;
    data[4107] =  'sd4244;
    data[4108] =  'sd21220;
    data[4109] = -'sd57741;
    data[4110] =  'sd38977;
    data[4111] =  'sd31044;
    data[4112] = -'sd8621;
    data[4113] = -'sd43105;
    data[4114] = -'sd51684;
    data[4115] =  'sd69262;
    data[4116] =  'sd18628;
    data[4117] = -'sd70701;
    data[4118] = -'sd25823;
    data[4119] =  'sd34726;
    data[4120] =  'sd9789;
    data[4121] =  'sd48945;
    data[4122] =  'sd80884;
    data[4123] =  'sd76738;
    data[4124] =  'sd56008;
    data[4125] = -'sd47642;
    data[4126] = -'sd74369;
    data[4127] = -'sd44163;
    data[4128] = -'sd56974;
    data[4129] =  'sd42812;
    data[4130] =  'sd50219;
    data[4131] = -'sd76587;
    data[4132] = -'sd55253;
    data[4133] =  'sd51417;
    data[4134] = -'sd70597;
    data[4135] = -'sd25303;
    data[4136] =  'sd37326;
    data[4137] =  'sd22789;
    data[4138] = -'sd49896;
    data[4139] =  'sd78202;
    data[4140] =  'sd63328;
    data[4141] = -'sd11042;
    data[4142] = -'sd55210;
    data[4143] =  'sd51632;
    data[4144] = -'sd69522;
    data[4145] = -'sd19928;
    data[4146] =  'sd64201;
    data[4147] = -'sd6677;
    data[4148] = -'sd33385;
    data[4149] = -'sd3084;
    data[4150] = -'sd15420;
    data[4151] = -'sd77100;
    data[4152] = -'sd57818;
    data[4153] =  'sd38592;
    data[4154] =  'sd29119;
    data[4155] = -'sd18246;
    data[4156] =  'sd72611;
    data[4157] =  'sd35373;
    data[4158] =  'sd13024;
    data[4159] =  'sd65120;
    data[4160] = -'sd2082;
    data[4161] = -'sd10410;
    data[4162] = -'sd52050;
    data[4163] =  'sd67432;
    data[4164] =  'sd9478;
    data[4165] =  'sd47390;
    data[4166] =  'sd73109;
    data[4167] =  'sd37863;
    data[4168] =  'sd25474;
    data[4169] = -'sd36471;
    data[4170] = -'sd18514;
    data[4171] =  'sd71271;
    data[4172] =  'sd28673;
    data[4173] = -'sd20476;
    data[4174] =  'sd61461;
    data[4175] = -'sd20377;
    data[4176] =  'sd61956;
    data[4177] = -'sd17902;
    data[4178] =  'sd74331;
    data[4179] =  'sd43973;
    data[4180] =  'sd56024;
    data[4181] = -'sd47562;
    data[4182] = -'sd73969;
    data[4183] = -'sd42163;
    data[4184] = -'sd46974;
    data[4185] = -'sd71029;
    data[4186] = -'sd27463;
    data[4187] =  'sd26526;
    data[4188] = -'sd31211;
    data[4189] =  'sd7786;
    data[4190] =  'sd38930;
    data[4191] =  'sd30809;
    data[4192] = -'sd9796;
    data[4193] = -'sd48980;
    data[4194] = -'sd81059;
    data[4195] = -'sd77613;
    data[4196] = -'sd60383;
    data[4197] =  'sd25767;
    data[4198] = -'sd35006;
    data[4199] = -'sd11189;
    data[4200] = -'sd55945;
    data[4201] =  'sd47957;
    data[4202] =  'sd75944;
    data[4203] =  'sd52038;
    data[4204] = -'sd67492;
    data[4205] = -'sd9778;
    data[4206] = -'sd48890;
    data[4207] = -'sd80609;
    data[4208] = -'sd75363;
    data[4209] = -'sd49133;
    data[4210] = -'sd81824;
    data[4211] = -'sd81438;
    data[4212] = -'sd79508;
    data[4213] = -'sd69858;
    data[4214] = -'sd21608;
    data[4215] =  'sd55801;
    data[4216] = -'sd48677;
    data[4217] = -'sd79544;
    data[4218] = -'sd70038;
    data[4219] = -'sd22508;
    data[4220] =  'sd51301;
    data[4221] = -'sd71177;
    data[4222] = -'sd28203;
    data[4223] =  'sd22826;
    data[4224] = -'sd49711;
    data[4225] =  'sd79127;
    data[4226] =  'sd67953;
    data[4227] =  'sd12083;
    data[4228] =  'sd60415;
    data[4229] = -'sd25607;
    data[4230] =  'sd35806;
    data[4231] =  'sd15189;
    data[4232] =  'sd75945;
    data[4233] =  'sd52043;
    data[4234] = -'sd67467;
    data[4235] = -'sd9653;
    data[4236] = -'sd48265;
    data[4237] = -'sd77484;
    data[4238] = -'sd59738;
    data[4239] =  'sd28992;
    data[4240] = -'sd18881;
    data[4241] =  'sd69436;
    data[4242] =  'sd19498;
    data[4243] = -'sd66351;
    data[4244] = -'sd4073;
    data[4245] = -'sd20365;
    data[4246] =  'sd62016;
    data[4247] = -'sd17602;
    data[4248] =  'sd75831;
    data[4249] =  'sd51473;
    data[4250] = -'sd70317;
    data[4251] = -'sd23903;
    data[4252] =  'sd44326;
    data[4253] =  'sd57789;
    data[4254] = -'sd38737;
    data[4255] = -'sd29844;
    data[4256] =  'sd14621;
    data[4257] =  'sd73105;
    data[4258] =  'sd37843;
    data[4259] =  'sd25374;
    data[4260] = -'sd36971;
    data[4261] = -'sd21014;
    data[4262] =  'sd58771;
    data[4263] = -'sd33827;
    data[4264] = -'sd5294;
    data[4265] = -'sd26470;
    data[4266] =  'sd31491;
    data[4267] = -'sd6386;
    data[4268] = -'sd31930;
    data[4269] =  'sd4191;
    data[4270] =  'sd20955;
    data[4271] = -'sd59066;
    data[4272] =  'sd32352;
    data[4273] = -'sd2081;
    data[4274] = -'sd10405;
    data[4275] = -'sd52025;
    data[4276] =  'sd67557;
    data[4277] =  'sd10103;
    data[4278] =  'sd50515;
    data[4279] = -'sd75107;
    data[4280] = -'sd47853;
    data[4281] = -'sd75424;
    data[4282] = -'sd49438;
    data[4283] =  'sd80492;
    data[4284] =  'sd74778;
    data[4285] =  'sd46208;
    data[4286] =  'sd67199;
    data[4287] =  'sd8313;
    data[4288] =  'sd41565;
    data[4289] =  'sd43984;
    data[4290] =  'sd56079;
    data[4291] = -'sd47287;
    data[4292] = -'sd72594;
    data[4293] = -'sd35288;
    data[4294] = -'sd12599;
    data[4295] = -'sd62995;
    data[4296] =  'sd12707;
    data[4297] =  'sd63535;
    data[4298] = -'sd10007;
    data[4299] = -'sd50035;
    data[4300] =  'sd77507;
    data[4301] =  'sd59853;
    data[4302] = -'sd28417;
    data[4303] =  'sd21756;
    data[4304] = -'sd55061;
    data[4305] =  'sd52377;
    data[4306] = -'sd65797;
    data[4307] = -'sd1303;
    data[4308] = -'sd6515;
    data[4309] = -'sd32575;
    data[4310] =  'sd966;
    data[4311] =  'sd4830;
    data[4312] =  'sd24150;
    data[4313] = -'sd43091;
    data[4314] = -'sd51614;
    data[4315] =  'sd69612;
    data[4316] =  'sd20378;
    data[4317] = -'sd61951;
    data[4318] =  'sd17927;
    data[4319] = -'sd74206;
    data[4320] = -'sd43348;
    data[4321] = -'sd52899;
    data[4322] =  'sd63187;
    data[4323] = -'sd11747;
    data[4324] = -'sd58735;
    data[4325] =  'sd34007;
    data[4326] =  'sd6194;
    data[4327] =  'sd30970;
    data[4328] = -'sd8991;
    data[4329] = -'sd44955;
    data[4330] = -'sd60934;
    data[4331] =  'sd23012;
    data[4332] = -'sd48781;
    data[4333] = -'sd80064;
    data[4334] = -'sd72638;
    data[4335] = -'sd35508;
    data[4336] = -'sd13699;
    data[4337] = -'sd68495;
    data[4338] = -'sd14793;
    data[4339] = -'sd73965;
    data[4340] = -'sd42143;
    data[4341] = -'sd46874;
    data[4342] = -'sd70529;
    data[4343] = -'sd24963;
    data[4344] =  'sd39026;
    data[4345] =  'sd31289;
    data[4346] = -'sd7396;
    data[4347] = -'sd36980;
    data[4348] = -'sd21059;
    data[4349] =  'sd58546;
    data[4350] = -'sd34952;
    data[4351] = -'sd10919;
    data[4352] = -'sd54595;
    data[4353] =  'sd54707;
    data[4354] = -'sd54147;
    data[4355] =  'sd56947;
    data[4356] = -'sd42947;
    data[4357] = -'sd50894;
    data[4358] =  'sd73212;
    data[4359] =  'sd38378;
    data[4360] =  'sd28049;
    data[4361] = -'sd23596;
    data[4362] =  'sd45861;
    data[4363] =  'sd65464;
    data[4364] = -'sd362;
    data[4365] = -'sd1810;
    data[4366] = -'sd9050;
    data[4367] = -'sd45250;
    data[4368] = -'sd62409;
    data[4369] =  'sd15637;
    data[4370] =  'sd78185;
    data[4371] =  'sd63243;
    data[4372] = -'sd11467;
    data[4373] = -'sd57335;
    data[4374] =  'sd41007;
    data[4375] =  'sd41194;
    data[4376] =  'sd42129;
    data[4377] =  'sd46804;
    data[4378] =  'sd70179;
    data[4379] =  'sd23213;
    data[4380] = -'sd47776;
    data[4381] = -'sd75039;
    data[4382] = -'sd47513;
    data[4383] = -'sd73724;
    data[4384] = -'sd40938;
    data[4385] = -'sd40849;
    data[4386] = -'sd40404;
    data[4387] = -'sd38179;
    data[4388] = -'sd27054;
    data[4389] =  'sd28571;
    data[4390] = -'sd20986;
    data[4391] =  'sd58911;
    data[4392] = -'sd33127;
    data[4393] = -'sd1794;
    data[4394] = -'sd8970;
    data[4395] = -'sd44850;
    data[4396] = -'sd60409;
    data[4397] =  'sd25637;
    data[4398] = -'sd35656;
    data[4399] = -'sd14439;
    data[4400] = -'sd72195;
    data[4401] = -'sd33293;
    data[4402] = -'sd2624;
    data[4403] = -'sd13120;
    data[4404] = -'sd65600;
    data[4405] = -'sd318;
    data[4406] = -'sd1590;
    data[4407] = -'sd7950;
    data[4408] = -'sd39750;
    data[4409] = -'sd34909;
    data[4410] = -'sd10704;
    data[4411] = -'sd53520;
    data[4412] =  'sd60082;
    data[4413] = -'sd27272;
    data[4414] =  'sd27481;
    data[4415] = -'sd26436;
    data[4416] =  'sd31661;
    data[4417] = -'sd5536;
    data[4418] = -'sd27680;
    data[4419] =  'sd25441;
    data[4420] = -'sd36636;
    data[4421] = -'sd19339;
    data[4422] =  'sd67146;
    data[4423] =  'sd8048;
    data[4424] =  'sd40240;
    data[4425] =  'sd37359;
    data[4426] =  'sd22954;
    data[4427] = -'sd49071;
    data[4428] = -'sd81514;
    data[4429] = -'sd79888;
    data[4430] = -'sd71758;
    data[4431] = -'sd31108;
    data[4432] =  'sd8301;
    data[4433] =  'sd41505;
    data[4434] =  'sd43684;
    data[4435] =  'sd54579;
    data[4436] = -'sd54787;
    data[4437] =  'sd53747;
    data[4438] = -'sd58947;
    data[4439] =  'sd32947;
    data[4440] =  'sd894;
    data[4441] =  'sd4470;
    data[4442] =  'sd22350;
    data[4443] = -'sd52091;
    data[4444] =  'sd67227;
    data[4445] =  'sd8453;
    data[4446] =  'sd42265;
    data[4447] =  'sd47484;
    data[4448] =  'sd73579;
    data[4449] =  'sd40213;
    data[4450] =  'sd37224;
    data[4451] =  'sd22279;
    data[4452] = -'sd52446;
    data[4453] =  'sd65452;
    data[4454] = -'sd422;
    data[4455] = -'sd2110;
    data[4456] = -'sd10550;
    data[4457] = -'sd52750;
    data[4458] =  'sd63932;
    data[4459] = -'sd8022;
    data[4460] = -'sd40110;
    data[4461] = -'sd36709;
    data[4462] = -'sd19704;
    data[4463] =  'sd65321;
    data[4464] = -'sd1077;
    data[4465] = -'sd5385;
    data[4466] = -'sd26925;
    data[4467] =  'sd29216;
    data[4468] = -'sd17761;
    data[4469] =  'sd75036;
    data[4470] =  'sd47498;
    data[4471] =  'sd73649;
    data[4472] =  'sd40563;
    data[4473] =  'sd38974;
    data[4474] =  'sd31029;
    data[4475] = -'sd8696;
    data[4476] = -'sd43480;
    data[4477] = -'sd53559;
    data[4478] =  'sd59887;
    data[4479] = -'sd28247;
    data[4480] =  'sd22606;
    data[4481] = -'sd50811;
    data[4482] =  'sd73627;
    data[4483] =  'sd40453;
    data[4484] =  'sd38424;
    data[4485] =  'sd28279;
    data[4486] = -'sd22446;
    data[4487] =  'sd51611;
    data[4488] = -'sd69627;
    data[4489] = -'sd20453;
    data[4490] =  'sd61576;
    data[4491] = -'sd19802;
    data[4492] =  'sd64831;
    data[4493] = -'sd3527;
    data[4494] = -'sd17635;
    data[4495] =  'sd75666;
    data[4496] =  'sd50648;
    data[4497] = -'sd74442;
    data[4498] = -'sd44528;
    data[4499] = -'sd58799;
    data[4500] =  'sd33687;
    data[4501] =  'sd4594;
    data[4502] =  'sd22970;
    data[4503] = -'sd48991;
    data[4504] = -'sd81114;
    data[4505] = -'sd77888;
    data[4506] = -'sd61758;
    data[4507] =  'sd18892;
    data[4508] = -'sd69381;
    data[4509] = -'sd19223;
    data[4510] =  'sd67726;
    data[4511] =  'sd10948;
    data[4512] =  'sd54740;
    data[4513] = -'sd53982;
    data[4514] =  'sd57772;
    data[4515] = -'sd38822;
    data[4516] = -'sd30269;
    data[4517] =  'sd12496;
    data[4518] =  'sd62480;
    data[4519] = -'sd15282;
    data[4520] = -'sd76410;
    data[4521] = -'sd54368;
    data[4522] =  'sd55842;
    data[4523] = -'sd48472;
    data[4524] = -'sd78519;
    data[4525] = -'sd64913;
    data[4526] =  'sd3117;
    data[4527] =  'sd15585;
    data[4528] =  'sd77925;
    data[4529] =  'sd61943;
    data[4530] = -'sd17967;
    data[4531] =  'sd74006;
    data[4532] =  'sd42348;
    data[4533] =  'sd47899;
    data[4534] =  'sd75654;
    data[4535] =  'sd50588;
    data[4536] = -'sd74742;
    data[4537] = -'sd46028;
    data[4538] = -'sd66299;
    data[4539] = -'sd3813;
    data[4540] = -'sd19065;
    data[4541] =  'sd68516;
    data[4542] =  'sd14898;
    data[4543] =  'sd74490;
    data[4544] =  'sd44768;
    data[4545] =  'sd59999;
    data[4546] = -'sd27687;
    data[4547] =  'sd25406;
    data[4548] = -'sd36811;
    data[4549] = -'sd20214;
    data[4550] =  'sd62771;
    data[4551] = -'sd13827;
    data[4552] = -'sd69135;
    data[4553] = -'sd17993;
    data[4554] =  'sd73876;
    data[4555] =  'sd41698;
    data[4556] =  'sd44649;
    data[4557] =  'sd59404;
    data[4558] = -'sd30662;
    data[4559] =  'sd10531;
    data[4560] =  'sd52655;
    data[4561] = -'sd64407;
    data[4562] =  'sd5647;
    data[4563] =  'sd28235;
    data[4564] = -'sd22666;
    data[4565] =  'sd50511;
    data[4566] = -'sd75127;
    data[4567] = -'sd47953;
    data[4568] = -'sd75924;
    data[4569] = -'sd51938;
    data[4570] =  'sd67992;
    data[4571] =  'sd12278;
    data[4572] =  'sd61390;
    data[4573] = -'sd20732;
    data[4574] =  'sd60181;
    data[4575] = -'sd26777;
    data[4576] =  'sd29956;
    data[4577] = -'sd14061;
    data[4578] = -'sd70305;
    data[4579] = -'sd23843;
    data[4580] =  'sd44626;
    data[4581] =  'sd59289;
    data[4582] = -'sd31237;
    data[4583] =  'sd7656;
    data[4584] =  'sd38280;
    data[4585] =  'sd27559;
    data[4586] = -'sd26046;
    data[4587] =  'sd33611;
    data[4588] =  'sd4214;
    data[4589] =  'sd21070;
    data[4590] = -'sd58491;
    data[4591] =  'sd35227;
    data[4592] =  'sd12294;
    data[4593] =  'sd61470;
    data[4594] = -'sd20332;
    data[4595] =  'sd62181;
    data[4596] = -'sd16777;
    data[4597] =  'sd79956;
    data[4598] =  'sd72098;
    data[4599] =  'sd32808;
    data[4600] =  'sd199;
    data[4601] =  'sd995;
    data[4602] =  'sd4975;
    data[4603] =  'sd24875;
    data[4604] = -'sd39466;
    data[4605] = -'sd33489;
    data[4606] = -'sd3604;
    data[4607] = -'sd18020;
    data[4608] =  'sd73741;
    data[4609] =  'sd41023;
    data[4610] =  'sd41274;
    data[4611] =  'sd42529;
    data[4612] =  'sd48804;
    data[4613] =  'sd80179;
    data[4614] =  'sd73213;
    data[4615] =  'sd38383;
    data[4616] =  'sd28074;
    data[4617] = -'sd23471;
    data[4618] =  'sd46486;
    data[4619] =  'sd68589;
    data[4620] =  'sd15263;
    data[4621] =  'sd76315;
    data[4622] =  'sd53893;
    data[4623] = -'sd58217;
    data[4624] =  'sd36597;
    data[4625] =  'sd19144;
    data[4626] = -'sd68121;
    data[4627] = -'sd12923;
    data[4628] = -'sd64615;
    data[4629] =  'sd4607;
    data[4630] =  'sd23035;
    data[4631] = -'sd48666;
    data[4632] = -'sd79489;
    data[4633] = -'sd69763;
    data[4634] = -'sd21133;
    data[4635] =  'sd58176;
    data[4636] = -'sd36802;
    data[4637] = -'sd20169;
    data[4638] =  'sd62996;
    data[4639] = -'sd12702;
    data[4640] = -'sd63510;
    data[4641] =  'sd10132;
    data[4642] =  'sd50660;
    data[4643] = -'sd74382;
    data[4644] = -'sd44228;
    data[4645] = -'sd57299;
    data[4646] =  'sd41187;
    data[4647] =  'sd42094;
    data[4648] =  'sd46629;
    data[4649] =  'sd69304;
    data[4650] =  'sd18838;
    data[4651] = -'sd69651;
    data[4652] = -'sd20573;
    data[4653] =  'sd60976;
    data[4654] = -'sd22802;
    data[4655] =  'sd49831;
    data[4656] = -'sd78527;
    data[4657] = -'sd64953;
    data[4658] =  'sd2917;
    data[4659] =  'sd14585;
    data[4660] =  'sd72925;
    data[4661] =  'sd36943;
    data[4662] =  'sd20874;
    data[4663] = -'sd59471;
    data[4664] =  'sd30327;
    data[4665] = -'sd12206;
    data[4666] = -'sd61030;
    data[4667] =  'sd22532;
    data[4668] = -'sd51181;
    data[4669] =  'sd71777;
    data[4670] =  'sd31203;
    data[4671] = -'sd7826;
    data[4672] = -'sd39130;
    data[4673] = -'sd31809;
    data[4674] =  'sd4796;
    data[4675] =  'sd23980;
    data[4676] = -'sd43941;
    data[4677] = -'sd55864;
    data[4678] =  'sd48362;
    data[4679] =  'sd77969;
    data[4680] =  'sd62163;
    data[4681] = -'sd16867;
    data[4682] =  'sd79506;
    data[4683] =  'sd69848;
    data[4684] =  'sd21558;
    data[4685] = -'sd56051;
    data[4686] =  'sd47427;
    data[4687] =  'sd73294;
    data[4688] =  'sd38788;
    data[4689] =  'sd30099;
    data[4690] = -'sd13346;
    data[4691] = -'sd66730;
    data[4692] = -'sd5968;
    data[4693] = -'sd29840;
    data[4694] =  'sd14641;
    data[4695] =  'sd73205;
    data[4696] =  'sd38343;
    data[4697] =  'sd27874;
    data[4698] = -'sd24471;
    data[4699] =  'sd41486;
    data[4700] =  'sd43589;
    data[4701] =  'sd54104;
    data[4702] = -'sd57162;
    data[4703] =  'sd41872;
    data[4704] =  'sd45519;
    data[4705] =  'sd63754;
    data[4706] = -'sd8912;
    data[4707] = -'sd44560;
    data[4708] = -'sd58959;
    data[4709] =  'sd32887;
    data[4710] =  'sd594;
    data[4711] =  'sd2970;
    data[4712] =  'sd14850;
    data[4713] =  'sd74250;
    data[4714] =  'sd43568;
    data[4715] =  'sd53999;
    data[4716] = -'sd57687;
    data[4717] =  'sd39247;
    data[4718] =  'sd32394;
    data[4719] = -'sd1871;
    data[4720] = -'sd9355;
    data[4721] = -'sd46775;
    data[4722] = -'sd70034;
    data[4723] = -'sd22488;
    data[4724] =  'sd51401;
    data[4725] = -'sd70677;
    data[4726] = -'sd25703;
    data[4727] =  'sd35326;
    data[4728] =  'sd12789;
    data[4729] =  'sd63945;
    data[4730] = -'sd7957;
    data[4731] = -'sd39785;
    data[4732] = -'sd35084;
    data[4733] = -'sd11579;
    data[4734] = -'sd57895;
    data[4735] =  'sd38207;
    data[4736] =  'sd27194;
    data[4737] = -'sd27871;
    data[4738] =  'sd24486;
    data[4739] = -'sd41411;
    data[4740] = -'sd43214;
    data[4741] = -'sd52229;
    data[4742] =  'sd66537;
    data[4743] =  'sd5003;
    data[4744] =  'sd25015;
    data[4745] = -'sd38766;
    data[4746] = -'sd29989;
    data[4747] =  'sd13896;
    data[4748] =  'sd69480;
    data[4749] =  'sd19718;
    data[4750] = -'sd65251;
    data[4751] =  'sd1427;
    data[4752] =  'sd7135;
    data[4753] =  'sd35675;
    data[4754] =  'sd14534;
    data[4755] =  'sd72670;
    data[4756] =  'sd35668;
    data[4757] =  'sd14499;
    data[4758] =  'sd72495;
    data[4759] =  'sd34793;
    data[4760] =  'sd10124;
    data[4761] =  'sd50620;
    data[4762] = -'sd74582;
    data[4763] = -'sd45228;
    data[4764] = -'sd62299;
    data[4765] =  'sd16187;
    data[4766] =  'sd80935;
    data[4767] =  'sd76993;
    data[4768] =  'sd57283;
    data[4769] = -'sd41267;
    data[4770] = -'sd42494;
    data[4771] = -'sd48629;
    data[4772] = -'sd79304;
    data[4773] = -'sd68838;
    data[4774] = -'sd16508;
    data[4775] =  'sd81301;
    data[4776] =  'sd78823;
    data[4777] =  'sd66433;
    data[4778] =  'sd4483;
    data[4779] =  'sd22415;
    data[4780] = -'sd51766;
    data[4781] =  'sd68852;
    data[4782] =  'sd16578;
    data[4783] = -'sd80951;
    data[4784] = -'sd77073;
    data[4785] = -'sd57683;
    data[4786] =  'sd39267;
    data[4787] =  'sd32494;
    data[4788] = -'sd1371;
    data[4789] = -'sd6855;
    data[4790] = -'sd34275;
    data[4791] = -'sd7534;
    data[4792] = -'sd37670;
    data[4793] = -'sd24509;
    data[4794] =  'sd41296;
    data[4795] =  'sd42639;
    data[4796] =  'sd49354;
    data[4797] = -'sd80912;
    data[4798] = -'sd76878;
    data[4799] = -'sd56708;
    data[4800] =  'sd44142;
    data[4801] =  'sd56869;
    data[4802] = -'sd43337;
    data[4803] = -'sd52844;
    data[4804] =  'sd63462;
    data[4805] = -'sd10372;
    data[4806] = -'sd51860;
    data[4807] =  'sd68382;
    data[4808] =  'sd14228;
    data[4809] =  'sd71140;
    data[4810] =  'sd28018;
    data[4811] = -'sd23751;
    data[4812] =  'sd45086;
    data[4813] =  'sd61589;
    data[4814] = -'sd19737;
    data[4815] =  'sd65156;
    data[4816] = -'sd1902;
    data[4817] = -'sd9510;
    data[4818] = -'sd47550;
    data[4819] = -'sd73909;
    data[4820] = -'sd41863;
    data[4821] = -'sd45474;
    data[4822] = -'sd63529;
    data[4823] =  'sd10037;
    data[4824] =  'sd50185;
    data[4825] = -'sd76757;
    data[4826] = -'sd56103;
    data[4827] =  'sd47167;
    data[4828] =  'sd71994;
    data[4829] =  'sd32288;
    data[4830] = -'sd2401;
    data[4831] = -'sd12005;
    data[4832] = -'sd60025;
    data[4833] =  'sd27557;
    data[4834] = -'sd26056;
    data[4835] =  'sd33561;
    data[4836] =  'sd3964;
    data[4837] =  'sd19820;
    data[4838] = -'sd64741;
    data[4839] =  'sd3977;
    data[4840] =  'sd19885;
    data[4841] = -'sd64416;
    data[4842] =  'sd5602;
    data[4843] =  'sd28010;
    data[4844] = -'sd23791;
    data[4845] =  'sd44886;
    data[4846] =  'sd60589;
    data[4847] = -'sd24737;
    data[4848] =  'sd40156;
    data[4849] =  'sd36939;
    data[4850] =  'sd20854;
    data[4851] = -'sd59571;
    data[4852] =  'sd29827;
    data[4853] = -'sd14706;
    data[4854] = -'sd73530;
    data[4855] = -'sd39968;
    data[4856] = -'sd35999;
    data[4857] = -'sd16154;
    data[4858] = -'sd80770;
    data[4859] = -'sd76168;
    data[4860] = -'sd53158;
    data[4861] =  'sd61892;
    data[4862] = -'sd18222;
    data[4863] =  'sd72731;
    data[4864] =  'sd35973;
    data[4865] =  'sd16024;
    data[4866] =  'sd80120;
    data[4867] =  'sd72918;
    data[4868] =  'sd36908;
    data[4869] =  'sd20699;
    data[4870] = -'sd60346;
    data[4871] =  'sd25952;
    data[4872] = -'sd34081;
    data[4873] = -'sd6564;
    data[4874] = -'sd32820;
    data[4875] = -'sd259;
    data[4876] = -'sd1295;
    data[4877] = -'sd6475;
    data[4878] = -'sd32375;
    data[4879] =  'sd1966;
    data[4880] =  'sd9830;
    data[4881] =  'sd49150;
    data[4882] =  'sd81909;
    data[4883] =  'sd81863;
    data[4884] =  'sd81633;
    data[4885] =  'sd80483;
    data[4886] =  'sd74733;
    data[4887] =  'sd45983;
    data[4888] =  'sd66074;
    data[4889] =  'sd2688;
    data[4890] =  'sd13440;
    data[4891] =  'sd67200;
    data[4892] =  'sd8318;
    data[4893] =  'sd41590;
    data[4894] =  'sd44109;
    data[4895] =  'sd56704;
    data[4896] = -'sd44162;
    data[4897] = -'sd56969;
    data[4898] =  'sd42837;
    data[4899] =  'sd50344;
    data[4900] = -'sd75962;
    data[4901] = -'sd52128;
    data[4902] =  'sd67042;
    data[4903] =  'sd7528;
    data[4904] =  'sd37640;
    data[4905] =  'sd24359;
    data[4906] = -'sd42046;
    data[4907] = -'sd46389;
    data[4908] = -'sd68104;
    data[4909] = -'sd12838;
    data[4910] = -'sd64190;
    data[4911] =  'sd6732;
    data[4912] =  'sd33660;
    data[4913] =  'sd4459;
    data[4914] =  'sd22295;
    data[4915] = -'sd52366;
    data[4916] =  'sd65852;
    data[4917] =  'sd1578;
    data[4918] =  'sd7890;
    data[4919] =  'sd39450;
    data[4920] =  'sd33409;
    data[4921] =  'sd3204;
    data[4922] =  'sd16020;
    data[4923] =  'sd80100;
    data[4924] =  'sd72818;
    data[4925] =  'sd36408;
    data[4926] =  'sd18199;
    data[4927] = -'sd72846;
    data[4928] = -'sd36548;
    data[4929] = -'sd18899;
    data[4930] =  'sd69346;
    data[4931] =  'sd19048;
    data[4932] = -'sd68601;
    data[4933] = -'sd15323;
    data[4934] = -'sd76615;
    data[4935] = -'sd55393;
    data[4936] =  'sd50717;
    data[4937] = -'sd74097;
    data[4938] = -'sd42803;
    data[4939] = -'sd50174;
    data[4940] =  'sd76812;
    data[4941] =  'sd56378;
    data[4942] = -'sd45792;
    data[4943] = -'sd65119;
    data[4944] =  'sd2087;
    data[4945] =  'sd10435;
    data[4946] =  'sd52175;
    data[4947] = -'sd66807;
    data[4948] = -'sd6353;
    data[4949] = -'sd31765;
    data[4950] =  'sd5016;
    data[4951] =  'sd25080;
    data[4952] = -'sd38441;
    data[4953] = -'sd28364;
    data[4954] =  'sd22021;
    data[4955] = -'sd53736;
    data[4956] =  'sd59002;
    data[4957] = -'sd32672;
    data[4958] =  'sd481;
    data[4959] =  'sd2405;
    data[4960] =  'sd12025;
    data[4961] =  'sd60125;
    data[4962] = -'sd27057;
    data[4963] =  'sd28556;
    data[4964] = -'sd21061;
    data[4965] =  'sd58536;
    data[4966] = -'sd35002;
    data[4967] = -'sd11169;
    data[4968] = -'sd55845;
    data[4969] =  'sd48457;
    data[4970] =  'sd78444;
    data[4971] =  'sd64538;
    data[4972] = -'sd4992;
    data[4973] = -'sd24960;
    data[4974] =  'sd39041;
    data[4975] =  'sd31364;
    data[4976] = -'sd7021;
    data[4977] = -'sd35105;
    data[4978] = -'sd11684;
    data[4979] = -'sd58420;
    data[4980] =  'sd35582;
    data[4981] =  'sd14069;
    data[4982] =  'sd70345;
    data[4983] =  'sd24043;
    data[4984] = -'sd43626;
    data[4985] = -'sd54289;
    data[4986] =  'sd56237;
    data[4987] = -'sd46497;
    data[4988] = -'sd68644;
    data[4989] = -'sd15538;
    data[4990] = -'sd77690;
    data[4991] = -'sd60768;
    data[4992] =  'sd23842;
    data[4993] = -'sd44631;
    data[4994] = -'sd59314;
    data[4995] =  'sd31112;
    data[4996] = -'sd8281;
    data[4997] = -'sd41405;
    data[4998] = -'sd43184;
    data[4999] = -'sd52079;
    data[5000] =  'sd67287;
    data[5001] =  'sd8753;
    data[5002] =  'sd43765;
    data[5003] =  'sd54984;
    data[5004] = -'sd52762;
    data[5005] =  'sd63872;
    data[5006] = -'sd8322;
    data[5007] = -'sd41610;
    data[5008] = -'sd44209;
    data[5009] = -'sd57204;
    data[5010] =  'sd41662;
    data[5011] =  'sd44469;
    data[5012] =  'sd58504;
    data[5013] = -'sd35162;
    data[5014] = -'sd11969;
    data[5015] = -'sd59845;
    data[5016] =  'sd28457;
    data[5017] = -'sd21556;
    data[5018] =  'sd56061;
    data[5019] = -'sd47377;
    data[5020] = -'sd73044;
    data[5021] = -'sd37538;
    data[5022] = -'sd23849;
    data[5023] =  'sd44596;
    data[5024] =  'sd59139;
    data[5025] = -'sd31987;
    data[5026] =  'sd3906;
    data[5027] =  'sd19530;
    data[5028] = -'sd66191;
    data[5029] = -'sd3273;
    data[5030] = -'sd16365;
    data[5031] = -'sd81825;
    data[5032] = -'sd81443;
    data[5033] = -'sd79533;
    data[5034] = -'sd69983;
    data[5035] = -'sd22233;
    data[5036] =  'sd52676;
    data[5037] = -'sd64302;
    data[5038] =  'sd6172;
    data[5039] =  'sd30860;
    data[5040] = -'sd9541;
    data[5041] = -'sd47705;
    data[5042] = -'sd74684;
    data[5043] = -'sd45738;
    data[5044] = -'sd64849;
    data[5045] =  'sd3437;
    data[5046] =  'sd17185;
    data[5047] = -'sd77916;
    data[5048] = -'sd61898;
    data[5049] =  'sd18192;
    data[5050] = -'sd72881;
    data[5051] = -'sd36723;
    data[5052] = -'sd19774;
    data[5053] =  'sd64971;
    data[5054] = -'sd2827;
    data[5055] = -'sd14135;
    data[5056] = -'sd70675;
    data[5057] = -'sd25693;
    data[5058] =  'sd35376;
    data[5059] =  'sd13039;
    data[5060] =  'sd65195;
    data[5061] = -'sd1707;
    data[5062] = -'sd8535;
    data[5063] = -'sd42675;
    data[5064] = -'sd49534;
    data[5065] =  'sd80012;
    data[5066] =  'sd72378;
    data[5067] =  'sd34208;
    data[5068] =  'sd7199;
    data[5069] =  'sd35995;
    data[5070] =  'sd16134;
    data[5071] =  'sd80670;
    data[5072] =  'sd75668;
    data[5073] =  'sd50658;
    data[5074] = -'sd74392;
    data[5075] = -'sd44278;
    data[5076] = -'sd57549;
    data[5077] =  'sd39937;
    data[5078] =  'sd35844;
    data[5079] =  'sd15379;
    data[5080] =  'sd76895;
    data[5081] =  'sd56793;
    data[5082] = -'sd43717;
    data[5083] = -'sd54744;
    data[5084] =  'sd53962;
    data[5085] = -'sd57872;
    data[5086] =  'sd38322;
    data[5087] =  'sd27769;
    data[5088] = -'sd24996;
    data[5089] =  'sd38861;
    data[5090] =  'sd30464;
    data[5091] = -'sd11521;
    data[5092] = -'sd57605;
    data[5093] =  'sd39657;
    data[5094] =  'sd34444;
    data[5095] =  'sd8379;
    data[5096] =  'sd41895;
    data[5097] =  'sd45634;
    data[5098] =  'sd64329;
    data[5099] = -'sd6037;
    data[5100] = -'sd30185;
    data[5101] =  'sd12916;
    data[5102] =  'sd64580;
    data[5103] = -'sd4782;
    data[5104] = -'sd23910;
    data[5105] =  'sd44291;
    data[5106] =  'sd57614;
    data[5107] = -'sd39612;
    data[5108] = -'sd34219;
    data[5109] = -'sd7254;
    data[5110] = -'sd36270;
    data[5111] = -'sd17509;
    data[5112] =  'sd76296;
    data[5113] =  'sd53798;
    data[5114] = -'sd58692;
    data[5115] =  'sd34222;
    data[5116] =  'sd7269;
    data[5117] =  'sd36345;
    data[5118] =  'sd17884;
    data[5119] = -'sd74421;
    data[5120] = -'sd44423;
    data[5121] = -'sd58274;
    data[5122] =  'sd36312;
    data[5123] =  'sd17719;
    data[5124] = -'sd75246;
    data[5125] = -'sd48548;
    data[5126] = -'sd78899;
    data[5127] = -'sd66813;
    data[5128] = -'sd6383;
    data[5129] = -'sd31915;
    data[5130] =  'sd4266;
    data[5131] =  'sd21330;
    data[5132] = -'sd57191;
    data[5133] =  'sd41727;
    data[5134] =  'sd44794;
    data[5135] =  'sd60129;
    data[5136] = -'sd27037;
    data[5137] =  'sd28656;
    data[5138] = -'sd20561;
    data[5139] =  'sd61036;
    data[5140] = -'sd22502;
    data[5141] =  'sd51331;
    data[5142] = -'sd71027;
    data[5143] = -'sd27453;
    data[5144] =  'sd26576;
    data[5145] = -'sd30961;
    data[5146] =  'sd9036;
    data[5147] =  'sd45180;
    data[5148] =  'sd62059;
    data[5149] = -'sd17387;
    data[5150] =  'sd76906;
    data[5151] =  'sd56848;
    data[5152] = -'sd43442;
    data[5153] = -'sd53369;
    data[5154] =  'sd60837;
    data[5155] = -'sd23497;
    data[5156] =  'sd46356;
    data[5157] =  'sd67939;
    data[5158] =  'sd12013;
    data[5159] =  'sd60065;
    data[5160] = -'sd27357;
    data[5161] =  'sd27056;
    data[5162] = -'sd28561;
    data[5163] =  'sd21036;
    data[5164] = -'sd58661;
    data[5165] =  'sd34377;
    data[5166] =  'sd8044;
    data[5167] =  'sd40220;
    data[5168] =  'sd37259;
    data[5169] =  'sd22454;
    data[5170] = -'sd51571;
    data[5171] =  'sd69827;
    data[5172] =  'sd21453;
    data[5173] = -'sd56576;
    data[5174] =  'sd44802;
    data[5175] =  'sd60169;
    data[5176] = -'sd26837;
    data[5177] =  'sd29656;
    data[5178] = -'sd15561;
    data[5179] = -'sd77805;
    data[5180] = -'sd61343;
    data[5181] =  'sd20967;
    data[5182] = -'sd59006;
    data[5183] =  'sd32652;
    data[5184] = -'sd581;
    data[5185] = -'sd2905;
    data[5186] = -'sd14525;
    data[5187] = -'sd72625;
    data[5188] = -'sd35443;
    data[5189] = -'sd13374;
    data[5190] = -'sd66870;
    data[5191] = -'sd6668;
    data[5192] = -'sd33340;
    data[5193] = -'sd2859;
    data[5194] = -'sd14295;
    data[5195] = -'sd71475;
    data[5196] = -'sd29693;
    data[5197] =  'sd15376;
    data[5198] =  'sd76880;
    data[5199] =  'sd56718;
    data[5200] = -'sd44092;
    data[5201] = -'sd56619;
    data[5202] =  'sd44587;
    data[5203] =  'sd59094;
    data[5204] = -'sd32212;
    data[5205] =  'sd2781;
    data[5206] =  'sd13905;
    data[5207] =  'sd69525;
    data[5208] =  'sd19943;
    data[5209] = -'sd64126;
    data[5210] =  'sd7052;
    data[5211] =  'sd35260;
    data[5212] =  'sd12459;
    data[5213] =  'sd62295;
    data[5214] = -'sd16207;
    data[5215] = -'sd81035;
    data[5216] = -'sd77493;
    data[5217] = -'sd59783;
    data[5218] =  'sd28767;
    data[5219] = -'sd20006;
    data[5220] =  'sd63811;
    data[5221] = -'sd8627;
    data[5222] = -'sd43135;
    data[5223] = -'sd51834;
    data[5224] =  'sd68512;
    data[5225] =  'sd14878;
    data[5226] =  'sd74390;
    data[5227] =  'sd44268;
    data[5228] =  'sd57499;
    data[5229] = -'sd40187;
    data[5230] = -'sd37094;
    data[5231] = -'sd21629;
    data[5232] =  'sd55696;
    data[5233] = -'sd49202;
    data[5234] =  'sd81672;
    data[5235] =  'sd80678;
    data[5236] =  'sd75708;
    data[5237] =  'sd50858;
    data[5238] = -'sd73392;
    data[5239] = -'sd39278;
    data[5240] = -'sd32549;
    data[5241] =  'sd1096;
    data[5242] =  'sd5480;
    data[5243] =  'sd27400;
    data[5244] = -'sd26841;
    data[5245] =  'sd29636;
    data[5246] = -'sd15661;
    data[5247] = -'sd78305;
    data[5248] = -'sd63843;
    data[5249] =  'sd8467;
    data[5250] =  'sd42335;
    data[5251] =  'sd47834;
    data[5252] =  'sd75329;
    data[5253] =  'sd48963;
    data[5254] =  'sd80974;
    data[5255] =  'sd77188;
    data[5256] =  'sd58258;
    data[5257] = -'sd36392;
    data[5258] = -'sd18119;
    data[5259] =  'sd73246;
    data[5260] =  'sd38548;
    data[5261] =  'sd28899;
    data[5262] = -'sd19346;
    data[5263] =  'sd67111;
    data[5264] =  'sd7873;
    data[5265] =  'sd39365;
    data[5266] =  'sd32984;
    data[5267] =  'sd1079;
    data[5268] =  'sd5395;
    data[5269] =  'sd26975;
    data[5270] = -'sd28966;
    data[5271] =  'sd19011;
    data[5272] = -'sd68786;
    data[5273] = -'sd16248;
    data[5274] = -'sd81240;
    data[5275] = -'sd78518;
    data[5276] = -'sd64908;
    data[5277] =  'sd3142;
    data[5278] =  'sd15710;
    data[5279] =  'sd78550;
    data[5280] =  'sd65068;
    data[5281] = -'sd2342;
    data[5282] = -'sd11710;
    data[5283] = -'sd58550;
    data[5284] =  'sd34932;
    data[5285] =  'sd10819;
    data[5286] =  'sd54095;
    data[5287] = -'sd57207;
    data[5288] =  'sd41647;
    data[5289] =  'sd44394;
    data[5290] =  'sd58129;
    data[5291] = -'sd37037;
    data[5292] = -'sd21344;
    data[5293] =  'sd57121;
    data[5294] = -'sd42077;
    data[5295] = -'sd46544;
    data[5296] = -'sd68879;
    data[5297] = -'sd16713;
    data[5298] =  'sd80276;
    data[5299] =  'sd73698;
    data[5300] =  'sd40808;
    data[5301] =  'sd40199;
    data[5302] =  'sd37154;
    data[5303] =  'sd21929;
    data[5304] = -'sd54196;
    data[5305] =  'sd56702;
    data[5306] = -'sd44172;
    data[5307] = -'sd57019;
    data[5308] =  'sd42587;
    data[5309] =  'sd49094;
    data[5310] =  'sd81629;
    data[5311] =  'sd80463;
    data[5312] =  'sd74633;
    data[5313] =  'sd45483;
    data[5314] =  'sd63574;
    data[5315] = -'sd9812;
    data[5316] = -'sd49060;
    data[5317] = -'sd81459;
    data[5318] = -'sd79613;
    data[5319] = -'sd70383;
    data[5320] = -'sd24233;
    data[5321] =  'sd42676;
    data[5322] =  'sd49539;
    data[5323] = -'sd79987;
    data[5324] = -'sd72253;
    data[5325] = -'sd33583;
    data[5326] = -'sd4074;
    data[5327] = -'sd20370;
    data[5328] =  'sd61991;
    data[5329] = -'sd17727;
    data[5330] =  'sd75206;
    data[5331] =  'sd48348;
    data[5332] =  'sd77899;
    data[5333] =  'sd61813;
    data[5334] = -'sd18617;
    data[5335] =  'sd70756;
    data[5336] =  'sd26098;
    data[5337] = -'sd33351;
    data[5338] = -'sd2914;
    data[5339] = -'sd14570;
    data[5340] = -'sd72850;
    data[5341] = -'sd36568;
    data[5342] = -'sd18999;
    data[5343] =  'sd68846;
    data[5344] =  'sd16548;
    data[5345] = -'sd81101;
    data[5346] = -'sd77823;
    data[5347] = -'sd61433;
    data[5348] =  'sd20517;
    data[5349] = -'sd61256;
    data[5350] =  'sd21402;
    data[5351] = -'sd56831;
    data[5352] =  'sd43527;
    data[5353] =  'sd53794;
    data[5354] = -'sd58712;
    data[5355] =  'sd34122;
    data[5356] =  'sd6769;
    data[5357] =  'sd33845;
    data[5358] =  'sd5384;
    data[5359] =  'sd26920;
    data[5360] = -'sd29241;
    data[5361] =  'sd17636;
    data[5362] = -'sd75661;
    data[5363] = -'sd50623;
    data[5364] =  'sd74567;
    data[5365] =  'sd45153;
    data[5366] =  'sd61924;
    data[5367] = -'sd18062;
    data[5368] =  'sd73531;
    data[5369] =  'sd39973;
    data[5370] =  'sd36024;
    data[5371] =  'sd16279;
    data[5372] =  'sd81395;
    data[5373] =  'sd79293;
    data[5374] =  'sd68783;
    data[5375] =  'sd16233;
    data[5376] =  'sd81165;
    data[5377] =  'sd78143;
    data[5378] =  'sd63033;
    data[5379] = -'sd12517;
    data[5380] = -'sd62585;
    data[5381] =  'sd14757;
    data[5382] =  'sd73785;
    data[5383] =  'sd41243;
    data[5384] =  'sd42374;
    data[5385] =  'sd48029;
    data[5386] =  'sd76304;
    data[5387] =  'sd53838;
    data[5388] = -'sd58492;
    data[5389] =  'sd35222;
    data[5390] =  'sd12269;
    data[5391] =  'sd61345;
    data[5392] = -'sd20957;
    data[5393] =  'sd59056;
    data[5394] = -'sd32402;
    data[5395] =  'sd1831;
    data[5396] =  'sd9155;
    data[5397] =  'sd45775;
    data[5398] =  'sd65034;
    data[5399] = -'sd2512;
    data[5400] = -'sd12560;
    data[5401] = -'sd62800;
    data[5402] =  'sd13682;
    data[5403] =  'sd68410;
    data[5404] =  'sd14368;
    data[5405] =  'sd71840;
    data[5406] =  'sd31518;
    data[5407] = -'sd6251;
    data[5408] = -'sd31255;
    data[5409] =  'sd7566;
    data[5410] =  'sd37830;
    data[5411] =  'sd25309;
    data[5412] = -'sd37296;
    data[5413] = -'sd22639;
    data[5414] =  'sd50646;
    data[5415] = -'sd74452;
    data[5416] = -'sd44578;
    data[5417] = -'sd59049;
    data[5418] =  'sd32437;
    data[5419] = -'sd1656;
    data[5420] = -'sd8280;
    data[5421] = -'sd41400;
    data[5422] = -'sd43159;
    data[5423] = -'sd51954;
    data[5424] =  'sd67912;
    data[5425] =  'sd11878;
    data[5426] =  'sd59390;
    data[5427] = -'sd30732;
    data[5428] =  'sd10181;
    data[5429] =  'sd50905;
    data[5430] = -'sd73157;
    data[5431] = -'sd38103;
    data[5432] = -'sd26674;
    data[5433] =  'sd30471;
    data[5434] = -'sd11486;
    data[5435] = -'sd57430;
    data[5436] =  'sd40532;
    data[5437] =  'sd38819;
    data[5438] =  'sd30254;
    data[5439] = -'sd12571;
    data[5440] = -'sd62855;
    data[5441] =  'sd13407;
    data[5442] =  'sd67035;
    data[5443] =  'sd7493;
    data[5444] =  'sd37465;
    data[5445] =  'sd23484;
    data[5446] = -'sd46421;
    data[5447] = -'sd68264;
    data[5448] = -'sd13638;
    data[5449] = -'sd68190;
    data[5450] = -'sd13268;
    data[5451] = -'sd66340;
    data[5452] = -'sd4018;
    data[5453] = -'sd20090;
    data[5454] =  'sd63391;
    data[5455] = -'sd10727;
    data[5456] = -'sd53635;
    data[5457] =  'sd59507;
    data[5458] = -'sd30147;
    data[5459] =  'sd13106;
    data[5460] =  'sd65530;
    data[5461] = -'sd32;
    data[5462] = -'sd160;
    data[5463] = -'sd800;
    data[5464] = -'sd4000;
    data[5465] = -'sd20000;
    data[5466] =  'sd63841;
    data[5467] = -'sd8477;
    data[5468] = -'sd42385;
    data[5469] = -'sd48084;
    data[5470] = -'sd76579;
    data[5471] = -'sd55213;
    data[5472] =  'sd51617;
    data[5473] = -'sd69597;
    data[5474] = -'sd20303;
    data[5475] =  'sd62326;
    data[5476] = -'sd16052;
    data[5477] = -'sd80260;
    data[5478] = -'sd73618;
    data[5479] = -'sd40408;
    data[5480] = -'sd38199;
    data[5481] = -'sd27154;
    data[5482] =  'sd28071;
    data[5483] = -'sd23486;
    data[5484] =  'sd46411;
    data[5485] =  'sd68214;
    data[5486] =  'sd13388;
    data[5487] =  'sd66940;
    data[5488] =  'sd7018;
    data[5489] =  'sd35090;
    data[5490] =  'sd11609;
    data[5491] =  'sd58045;
    data[5492] = -'sd37457;
    data[5493] = -'sd23444;
    data[5494] =  'sd46621;
    data[5495] =  'sd69264;
    data[5496] =  'sd18638;
    data[5497] = -'sd70651;
    data[5498] = -'sd25573;
    data[5499] =  'sd35976;
    data[5500] =  'sd16039;
    data[5501] =  'sd80195;
    data[5502] =  'sd73293;
    data[5503] =  'sd38783;
    data[5504] =  'sd30074;
    data[5505] = -'sd13471;
    data[5506] = -'sd67355;
    data[5507] = -'sd9093;
    data[5508] = -'sd45465;
    data[5509] = -'sd63484;
    data[5510] =  'sd10262;
    data[5511] =  'sd51310;
    data[5512] = -'sd71132;
    data[5513] = -'sd27978;
    data[5514] =  'sd23951;
    data[5515] = -'sd44086;
    data[5516] = -'sd56589;
    data[5517] =  'sd44737;
    data[5518] =  'sd59844;
    data[5519] = -'sd28462;
    data[5520] =  'sd21531;
    data[5521] = -'sd56186;
    data[5522] =  'sd46752;
    data[5523] =  'sd69919;
    data[5524] =  'sd21913;
    data[5525] = -'sd54276;
    data[5526] =  'sd56302;
    data[5527] = -'sd46172;
    data[5528] = -'sd67019;
    data[5529] = -'sd7413;
    data[5530] = -'sd37065;
    data[5531] = -'sd21484;
    data[5532] =  'sd56421;
    data[5533] = -'sd45577;
    data[5534] = -'sd64044;
    data[5535] =  'sd7462;
    data[5536] =  'sd37310;
    data[5537] =  'sd22709;
    data[5538] = -'sd50296;
    data[5539] =  'sd76202;
    data[5540] =  'sd53328;
    data[5541] = -'sd61042;
    data[5542] =  'sd22472;
    data[5543] = -'sd51481;
    data[5544] =  'sd70277;
    data[5545] =  'sd23703;
    data[5546] = -'sd45326;
    data[5547] = -'sd62789;
    data[5548] =  'sd13737;
    data[5549] =  'sd68685;
    data[5550] =  'sd15743;
    data[5551] =  'sd78715;
    data[5552] =  'sd65893;
    data[5553] =  'sd1783;
    data[5554] =  'sd8915;
    data[5555] =  'sd44575;
    data[5556] =  'sd59034;
    data[5557] = -'sd32512;
    data[5558] =  'sd1281;
    data[5559] =  'sd6405;
    data[5560] =  'sd32025;
    data[5561] = -'sd3716;
    data[5562] = -'sd18580;
    data[5563] =  'sd70941;
    data[5564] =  'sd27023;
    data[5565] = -'sd28726;
    data[5566] =  'sd20211;
    data[5567] = -'sd62786;
    data[5568] =  'sd13752;
    data[5569] =  'sd68760;
    data[5570] =  'sd16118;
    data[5571] =  'sd80590;
    data[5572] =  'sd75268;
    data[5573] =  'sd48658;
    data[5574] =  'sd79449;
    data[5575] =  'sd69563;
    data[5576] =  'sd20133;
    data[5577] = -'sd63176;
    data[5578] =  'sd11802;
    data[5579] =  'sd59010;
    data[5580] = -'sd32632;
    data[5581] =  'sd681;
    data[5582] =  'sd3405;
    data[5583] =  'sd17025;
    data[5584] = -'sd78716;
    data[5585] = -'sd65898;
    data[5586] = -'sd1808;
    data[5587] = -'sd9040;
    data[5588] = -'sd45200;
    data[5589] = -'sd62159;
    data[5590] =  'sd16887;
    data[5591] = -'sd79406;
    data[5592] = -'sd69348;
    data[5593] = -'sd19058;
    data[5594] =  'sd68551;
    data[5595] =  'sd15073;
    data[5596] =  'sd75365;
    data[5597] =  'sd49143;
    data[5598] =  'sd81874;
    data[5599] =  'sd81688;
    data[5600] =  'sd80758;
    data[5601] =  'sd76108;
    data[5602] =  'sd52858;
    data[5603] = -'sd63392;
    data[5604] =  'sd10722;
    data[5605] =  'sd53610;
    data[5606] = -'sd59632;
    data[5607] =  'sd29522;
    data[5608] = -'sd16231;
    data[5609] = -'sd81155;
    data[5610] = -'sd78093;
    data[5611] = -'sd62783;
    data[5612] =  'sd13767;
    data[5613] =  'sd68835;
    data[5614] =  'sd16493;
    data[5615] = -'sd81376;
    data[5616] = -'sd79198;
    data[5617] = -'sd68308;
    data[5618] = -'sd13858;
    data[5619] = -'sd69290;
    data[5620] = -'sd18768;
    data[5621] =  'sd70001;
    data[5622] =  'sd22323;
    data[5623] = -'sd52226;
    data[5624] =  'sd66552;
    data[5625] =  'sd5078;
    data[5626] =  'sd25390;
    data[5627] = -'sd36891;
    data[5628] = -'sd20614;
    data[5629] =  'sd60771;
    data[5630] = -'sd23827;
    data[5631] =  'sd44706;
    data[5632] =  'sd59689;
    data[5633] = -'sd29237;
    data[5634] =  'sd17656;
    data[5635] = -'sd75561;
    data[5636] = -'sd50123;
    data[5637] =  'sd77067;
    data[5638] =  'sd57653;
    data[5639] = -'sd39417;
    data[5640] = -'sd33244;
    data[5641] = -'sd2379;
    data[5642] = -'sd11895;
    data[5643] = -'sd59475;
    data[5644] =  'sd30307;
    data[5645] = -'sd12306;
    data[5646] = -'sd61530;
    data[5647] =  'sd20032;
    data[5648] = -'sd63681;
    data[5649] =  'sd9277;
    data[5650] =  'sd46385;
    data[5651] =  'sd68084;
    data[5652] =  'sd12738;
    data[5653] =  'sd63690;
    data[5654] = -'sd9232;
    data[5655] = -'sd46160;
    data[5656] = -'sd66959;
    data[5657] = -'sd7113;
    data[5658] = -'sd35565;
    data[5659] = -'sd13984;
    data[5660] = -'sd69920;
    data[5661] = -'sd21918;
    data[5662] =  'sd54251;
    data[5663] = -'sd56427;
    data[5664] =  'sd45547;
    data[5665] =  'sd63894;
    data[5666] = -'sd8212;
    data[5667] = -'sd41060;
    data[5668] = -'sd41459;
    data[5669] = -'sd43454;
    data[5670] = -'sd53429;
    data[5671] =  'sd60537;
    data[5672] = -'sd24997;
    data[5673] =  'sd38856;
    data[5674] =  'sd30439;
    data[5675] = -'sd11646;
    data[5676] = -'sd58230;
    data[5677] =  'sd36532;
    data[5678] =  'sd18819;
    data[5679] = -'sd69746;
    data[5680] = -'sd21048;
    data[5681] =  'sd58601;
    data[5682] = -'sd34677;
    data[5683] = -'sd9544;
    data[5684] = -'sd47720;
    data[5685] = -'sd74759;
    data[5686] = -'sd46113;
    data[5687] = -'sd66724;
    data[5688] = -'sd5938;
    data[5689] = -'sd29690;
    data[5690] =  'sd15391;
    data[5691] =  'sd76955;
    data[5692] =  'sd57093;
    data[5693] = -'sd42217;
    data[5694] = -'sd47244;
    data[5695] = -'sd72379;
    data[5696] = -'sd34213;
    data[5697] = -'sd7224;
    data[5698] = -'sd36120;
    data[5699] = -'sd16759;
    data[5700] =  'sd80046;
    data[5701] =  'sd72548;
    data[5702] =  'sd35058;
    data[5703] =  'sd11449;
    data[5704] =  'sd57245;
    data[5705] = -'sd41457;
    data[5706] = -'sd43444;
    data[5707] = -'sd53379;
    data[5708] =  'sd60787;
    data[5709] = -'sd23747;
    data[5710] =  'sd45106;
    data[5711] =  'sd61689;
    data[5712] = -'sd19237;
    data[5713] =  'sd67656;
    data[5714] =  'sd10598;
    data[5715] =  'sd52990;
    data[5716] = -'sd62732;
    data[5717] =  'sd14022;
    data[5718] =  'sd70110;
    data[5719] =  'sd22868;
    data[5720] = -'sd49501;
    data[5721] =  'sd80177;
    data[5722] =  'sd73203;
    data[5723] =  'sd38333;
    data[5724] =  'sd27824;
    data[5725] = -'sd24721;
    data[5726] =  'sd40236;
    data[5727] =  'sd37339;
    data[5728] =  'sd22854;
    data[5729] = -'sd49571;
    data[5730] =  'sd79827;
    data[5731] =  'sd71453;
    data[5732] =  'sd29583;
    data[5733] = -'sd15926;
    data[5734] = -'sd79630;
    data[5735] = -'sd70468;
    data[5736] = -'sd24658;
    data[5737] =  'sd40551;
    data[5738] =  'sd38914;
    data[5739] =  'sd30729;
    data[5740] = -'sd10196;
    data[5741] = -'sd50980;
    data[5742] =  'sd72782;
    data[5743] =  'sd36228;
    data[5744] =  'sd17299;
    data[5745] = -'sd77346;
    data[5746] = -'sd59048;
    data[5747] =  'sd32442;
    data[5748] = -'sd1631;
    data[5749] = -'sd8155;
    data[5750] = -'sd40775;
    data[5751] = -'sd40034;
    data[5752] = -'sd36329;
    data[5753] = -'sd17804;
    data[5754] =  'sd74821;
    data[5755] =  'sd46423;
    data[5756] =  'sd68274;
    data[5757] =  'sd13688;
    data[5758] =  'sd68440;
    data[5759] =  'sd14518;
    data[5760] =  'sd72590;
    data[5761] =  'sd35268;
    data[5762] =  'sd12499;
    data[5763] =  'sd62495;
    data[5764] = -'sd15207;
    data[5765] = -'sd76035;
    data[5766] = -'sd52493;
    data[5767] =  'sd65217;
    data[5768] = -'sd1597;
    data[5769] = -'sd7985;
    data[5770] = -'sd39925;
    data[5771] = -'sd35784;
    data[5772] = -'sd15079;
    data[5773] = -'sd75395;
    data[5774] = -'sd49293;
    data[5775] =  'sd81217;
    data[5776] =  'sd78403;
    data[5777] =  'sd64333;
    data[5778] = -'sd6017;
    data[5779] = -'sd30085;
    data[5780] =  'sd13416;
    data[5781] =  'sd67080;
    data[5782] =  'sd7718;
    data[5783] =  'sd38590;
    data[5784] =  'sd29109;
    data[5785] = -'sd18296;
    data[5786] =  'sd72361;
    data[5787] =  'sd34123;
    data[5788] =  'sd6774;
    data[5789] =  'sd33870;
    data[5790] =  'sd5509;
    data[5791] =  'sd27545;
    data[5792] = -'sd26116;
    data[5793] =  'sd33261;
    data[5794] =  'sd2464;
    data[5795] =  'sd12320;
    data[5796] =  'sd61600;
    data[5797] = -'sd19682;
    data[5798] =  'sd65431;
    data[5799] = -'sd527;
    data[5800] = -'sd2635;
    data[5801] = -'sd13175;
    data[5802] = -'sd65875;
    data[5803] = -'sd1693;
    data[5804] = -'sd8465;
    data[5805] = -'sd42325;
    data[5806] = -'sd47784;
    data[5807] = -'sd75079;
    data[5808] = -'sd47713;
    data[5809] = -'sd74724;
    data[5810] = -'sd45938;
    data[5811] = -'sd65849;
    data[5812] = -'sd1563;
    data[5813] = -'sd7815;
    data[5814] = -'sd39075;
    data[5815] = -'sd31534;
    data[5816] =  'sd6171;
    data[5817] =  'sd30855;
    data[5818] = -'sd9566;
    data[5819] = -'sd47830;
    data[5820] = -'sd75309;
    data[5821] = -'sd48863;
    data[5822] = -'sd80474;
    data[5823] = -'sd74688;
    data[5824] = -'sd45758;
    data[5825] = -'sd64949;
    data[5826] =  'sd2937;
    data[5827] =  'sd14685;
    data[5828] =  'sd73425;
    data[5829] =  'sd39443;
    data[5830] =  'sd33374;
    data[5831] =  'sd3029;
    data[5832] =  'sd15145;
    data[5833] =  'sd75725;
    data[5834] =  'sd50943;
    data[5835] = -'sd72967;
    data[5836] = -'sd37153;
    data[5837] = -'sd21924;
    data[5838] =  'sd54221;
    data[5839] = -'sd56577;
    data[5840] =  'sd44797;
    data[5841] =  'sd60144;
    data[5842] = -'sd26962;
    data[5843] =  'sd29031;
    data[5844] = -'sd18686;
    data[5845] =  'sd70411;
    data[5846] =  'sd24373;
    data[5847] = -'sd41976;
    data[5848] = -'sd46039;
    data[5849] = -'sd66354;
    data[5850] = -'sd4088;
    data[5851] = -'sd20440;
    data[5852] =  'sd61641;
    data[5853] = -'sd19477;
    data[5854] =  'sd66456;
    data[5855] =  'sd4598;
    data[5856] =  'sd22990;
    data[5857] = -'sd48891;
    data[5858] = -'sd80614;
    data[5859] = -'sd75388;
    data[5860] = -'sd49258;
    data[5861] =  'sd81392;
    data[5862] =  'sd79278;
    data[5863] =  'sd68708;
    data[5864] =  'sd15858;
    data[5865] =  'sd79290;
    data[5866] =  'sd68768;
    data[5867] =  'sd16158;
    data[5868] =  'sd80790;
    data[5869] =  'sd76268;
    data[5870] =  'sd53658;
    data[5871] = -'sd59392;
    data[5872] =  'sd30722;
    data[5873] = -'sd10231;
    data[5874] = -'sd51155;
    data[5875] =  'sd71907;
    data[5876] =  'sd31853;
    data[5877] = -'sd4576;
    data[5878] = -'sd22880;
    data[5879] =  'sd49441;
    data[5880] = -'sd80477;
    data[5881] = -'sd74703;
    data[5882] = -'sd45833;
    data[5883] = -'sd65324;
    data[5884] =  'sd1062;
    data[5885] =  'sd5310;
    data[5886] =  'sd26550;
    data[5887] = -'sd31091;
    data[5888] =  'sd8386;
    data[5889] =  'sd41930;
    data[5890] =  'sd45809;
    data[5891] =  'sd65204;
    data[5892] = -'sd1662;
    data[5893] = -'sd8310;
    data[5894] = -'sd41550;
    data[5895] = -'sd43909;
    data[5896] = -'sd55704;
    data[5897] =  'sd49162;
    data[5898] = -'sd81872;
    data[5899] = -'sd81678;
    data[5900] = -'sd80708;
    data[5901] = -'sd75858;
    data[5902] = -'sd51608;
    data[5903] =  'sd69642;
    data[5904] =  'sd20528;
    data[5905] = -'sd61201;
    data[5906] =  'sd21677;
    data[5907] = -'sd55456;
    data[5908] =  'sd50402;
    data[5909] = -'sd75672;
    data[5910] = -'sd50678;
    data[5911] =  'sd74292;
    data[5912] =  'sd43778;
    data[5913] =  'sd55049;
    data[5914] = -'sd52437;
    data[5915] =  'sd65497;
    data[5916] = -'sd197;
    data[5917] = -'sd985;
    data[5918] = -'sd4925;
    data[5919] = -'sd24625;
    data[5920] =  'sd40716;
    data[5921] =  'sd39739;
    data[5922] =  'sd34854;
    data[5923] =  'sd10429;
    data[5924] =  'sd52145;
    data[5925] = -'sd66957;
    data[5926] = -'sd7103;
    data[5927] = -'sd35515;
    data[5928] = -'sd13734;
    data[5929] = -'sd68670;
    data[5930] = -'sd15668;
    data[5931] = -'sd78340;
    data[5932] = -'sd64018;
    data[5933] =  'sd7592;
    data[5934] =  'sd37960;
    data[5935] =  'sd25959;
    data[5936] = -'sd34046;
    data[5937] = -'sd6389;
    data[5938] = -'sd31945;
    data[5939] =  'sd4116;
    data[5940] =  'sd20580;
    data[5941] = -'sd60941;
    data[5942] =  'sd22977;
    data[5943] = -'sd48956;
    data[5944] = -'sd80939;
    data[5945] = -'sd77013;
    data[5946] = -'sd57383;
    data[5947] =  'sd40767;
    data[5948] =  'sd39994;
    data[5949] =  'sd36129;
    data[5950] =  'sd16804;
    data[5951] = -'sd79821;
    data[5952] = -'sd71423;
    data[5953] = -'sd29433;
    data[5954] =  'sd16676;
    data[5955] = -'sd80461;
    data[5956] = -'sd74623;
    data[5957] = -'sd45433;
    data[5958] = -'sd63324;
    data[5959] =  'sd11062;
    data[5960] =  'sd55310;
    data[5961] = -'sd51132;
    data[5962] =  'sd72022;
    data[5963] =  'sd32428;
    data[5964] = -'sd1701;
    data[5965] = -'sd8505;
    data[5966] = -'sd42525;
    data[5967] = -'sd48784;
    data[5968] = -'sd80079;
    data[5969] = -'sd72713;
    data[5970] = -'sd35883;
    data[5971] = -'sd15574;
    data[5972] = -'sd77870;
    data[5973] = -'sd61668;
    data[5974] =  'sd19342;
    data[5975] = -'sd67131;
    data[5976] = -'sd7973;
    data[5977] = -'sd39865;
    data[5978] = -'sd35484;
    data[5979] = -'sd13579;
    data[5980] = -'sd67895;
    data[5981] = -'sd11793;
    data[5982] = -'sd58965;
    data[5983] =  'sd32857;
    data[5984] =  'sd444;
    data[5985] =  'sd2220;
    data[5986] =  'sd11100;
    data[5987] =  'sd55500;
    data[5988] = -'sd50182;
    data[5989] =  'sd76772;
    data[5990] =  'sd56178;
    data[5991] = -'sd46792;
    data[5992] = -'sd70119;
    data[5993] = -'sd22913;
    data[5994] =  'sd49276;
    data[5995] = -'sd81302;
    data[5996] = -'sd78828;
    data[5997] = -'sd66458;
    data[5998] = -'sd4608;
    data[5999] = -'sd23040;
    data[6000] =  'sd48641;
    data[6001] =  'sd79364;
    data[6002] =  'sd69138;
    data[6003] =  'sd18008;
    data[6004] = -'sd73801;
    data[6005] = -'sd41323;
    data[6006] = -'sd42774;
    data[6007] = -'sd50029;
    data[6008] =  'sd77537;
    data[6009] =  'sd60003;
    data[6010] = -'sd27667;
    data[6011] =  'sd25506;
    data[6012] = -'sd36311;
    data[6013] = -'sd17714;
    data[6014] =  'sd75271;
    data[6015] =  'sd48673;
    data[6016] =  'sd79524;
    data[6017] =  'sd69938;
    data[6018] =  'sd22008;
    data[6019] = -'sd53801;
    data[6020] =  'sd58677;
    data[6021] = -'sd34297;
    data[6022] = -'sd7644;
    data[6023] = -'sd38220;
    data[6024] = -'sd27259;
    data[6025] =  'sd27546;
    data[6026] = -'sd26111;
    data[6027] =  'sd33286;
    data[6028] =  'sd2589;
    data[6029] =  'sd12945;
    data[6030] =  'sd64725;
    data[6031] = -'sd4057;
    data[6032] = -'sd20285;
    data[6033] =  'sd62416;
    data[6034] = -'sd15602;
    data[6035] = -'sd78010;
    data[6036] = -'sd62368;
    data[6037] =  'sd15842;
    data[6038] =  'sd79210;
    data[6039] =  'sd68368;
    data[6040] =  'sd14158;
    data[6041] =  'sd70790;
    data[6042] =  'sd26268;
    data[6043] = -'sd32501;
    data[6044] =  'sd1336;
    data[6045] =  'sd6680;
    data[6046] =  'sd33400;
    data[6047] =  'sd3159;
    data[6048] =  'sd15795;
    data[6049] =  'sd78975;
    data[6050] =  'sd67193;
    data[6051] =  'sd8283;
    data[6052] =  'sd41415;
    data[6053] =  'sd43234;
    data[6054] =  'sd52329;
    data[6055] = -'sd66037;
    data[6056] = -'sd2503;
    data[6057] = -'sd12515;
    data[6058] = -'sd62575;
    data[6059] =  'sd14807;
    data[6060] =  'sd74035;
    data[6061] =  'sd42493;
    data[6062] =  'sd48624;
    data[6063] =  'sd79279;
    data[6064] =  'sd68713;
    data[6065] =  'sd15883;
    data[6066] =  'sd79415;
    data[6067] =  'sd69393;
    data[6068] =  'sd19283;
    data[6069] = -'sd67426;
    data[6070] = -'sd9448;
    data[6071] = -'sd47240;
    data[6072] = -'sd72359;
    data[6073] = -'sd34113;
    data[6074] = -'sd6724;
    data[6075] = -'sd33620;
    data[6076] = -'sd4259;
    data[6077] = -'sd21295;
    data[6078] =  'sd57366;
    data[6079] = -'sd40852;
    data[6080] = -'sd40419;
    data[6081] = -'sd38254;
    data[6082] = -'sd27429;
    data[6083] =  'sd26696;
    data[6084] = -'sd30361;
    data[6085] =  'sd12036;
    data[6086] =  'sd60180;
    data[6087] = -'sd26782;
    data[6088] =  'sd29931;
    data[6089] = -'sd14186;
    data[6090] = -'sd70930;
    data[6091] = -'sd26968;
    data[6092] =  'sd29001;
    data[6093] = -'sd18836;
    data[6094] =  'sd69661;
    data[6095] =  'sd20623;
    data[6096] = -'sd60726;
    data[6097] =  'sd24052;
    data[6098] = -'sd43581;
    data[6099] = -'sd54064;
    data[6100] =  'sd57362;
    data[6101] = -'sd40872;
    data[6102] = -'sd40519;
    data[6103] = -'sd38754;
    data[6104] = -'sd29929;
    data[6105] =  'sd14196;
    data[6106] =  'sd70980;
    data[6107] =  'sd27218;
    data[6108] = -'sd27751;
    data[6109] =  'sd25086;
    data[6110] = -'sd38411;
    data[6111] = -'sd28214;
    data[6112] =  'sd22771;
    data[6113] = -'sd49986;
    data[6114] =  'sd77752;
    data[6115] =  'sd61078;
    data[6116] = -'sd22292;
    data[6117] =  'sd52381;
    data[6118] = -'sd65777;
    data[6119] = -'sd1203;
    data[6120] = -'sd6015;
    data[6121] = -'sd30075;
    data[6122] =  'sd13466;
    data[6123] =  'sd67330;
    data[6124] =  'sd8968;
    data[6125] =  'sd44840;
    data[6126] =  'sd60359;
    data[6127] = -'sd25887;
    data[6128] =  'sd34406;
    data[6129] =  'sd8189;
    data[6130] =  'sd40945;
    data[6131] =  'sd40884;
    data[6132] =  'sd40579;
    data[6133] =  'sd39054;
    data[6134] =  'sd31429;
    data[6135] = -'sd6696;
    data[6136] = -'sd33480;
    data[6137] = -'sd3559;
    data[6138] = -'sd17795;
    data[6139] =  'sd74866;
    data[6140] =  'sd46648;
    data[6141] =  'sd69399;
    data[6142] =  'sd19313;
    data[6143] = -'sd67276;
    data[6144] = -'sd8698;
    data[6145] = -'sd43490;
    data[6146] = -'sd53609;
    data[6147] =  'sd59637;
    data[6148] = -'sd29497;
    data[6149] =  'sd16356;
    data[6150] =  'sd81780;
    data[6151] =  'sd81218;
    data[6152] =  'sd78408;
    data[6153] =  'sd64358;
    data[6154] = -'sd5892;
    data[6155] = -'sd29460;
    data[6156] =  'sd16541;
    data[6157] = -'sd81136;
    data[6158] = -'sd77998;
    data[6159] = -'sd62308;
    data[6160] =  'sd16142;
    data[6161] =  'sd80710;
    data[6162] =  'sd75868;
    data[6163] =  'sd51658;
    data[6164] = -'sd69392;
    data[6165] = -'sd19278;
    data[6166] =  'sd67451;
    data[6167] =  'sd9573;
    data[6168] =  'sd47865;
    data[6169] =  'sd75484;
    data[6170] =  'sd49738;
    data[6171] = -'sd78992;
    data[6172] = -'sd67278;
    data[6173] = -'sd8708;
    data[6174] = -'sd43540;
    data[6175] = -'sd53859;
    data[6176] =  'sd58387;
    data[6177] = -'sd35747;
    data[6178] = -'sd14894;
    data[6179] = -'sd74470;
    data[6180] = -'sd44668;
    data[6181] = -'sd59499;
    data[6182] =  'sd30187;
    data[6183] = -'sd12906;
    data[6184] = -'sd64530;
    data[6185] =  'sd5032;
    data[6186] =  'sd25160;
    data[6187] = -'sd38041;
    data[6188] = -'sd26364;
    data[6189] =  'sd32021;
    data[6190] = -'sd3736;
    data[6191] = -'sd18680;
    data[6192] =  'sd70441;
    data[6193] =  'sd24523;
    data[6194] = -'sd41226;
    data[6195] = -'sd42289;
    data[6196] = -'sd47604;
    data[6197] = -'sd74179;
    data[6198] = -'sd43213;
    data[6199] = -'sd52224;
    data[6200] =  'sd66562;
    data[6201] =  'sd5128;
    data[6202] =  'sd25640;
    data[6203] = -'sd35641;
    data[6204] = -'sd14364;
    data[6205] = -'sd71820;
    data[6206] = -'sd31418;
    data[6207] =  'sd6751;
    data[6208] =  'sd33755;
    data[6209] =  'sd4934;
    data[6210] =  'sd24670;
    data[6211] = -'sd40491;
    data[6212] = -'sd38614;
    data[6213] = -'sd29229;
    data[6214] =  'sd17696;
    data[6215] = -'sd75361;
    data[6216] = -'sd49123;
    data[6217] = -'sd81774;
    data[6218] = -'sd81188;
    data[6219] = -'sd78258;
    data[6220] = -'sd63608;
    data[6221] =  'sd9642;
    data[6222] =  'sd48210;
    data[6223] =  'sd77209;
    data[6224] =  'sd58363;
    data[6225] = -'sd35867;
    data[6226] = -'sd15494;
    data[6227] = -'sd77470;
    data[6228] = -'sd59668;
    data[6229] =  'sd29342;
    data[6230] = -'sd17131;
    data[6231] =  'sd78186;
    data[6232] =  'sd63248;
    data[6233] = -'sd11442;
    data[6234] = -'sd57210;
    data[6235] =  'sd41632;
    data[6236] =  'sd44319;
    data[6237] =  'sd57754;
    data[6238] = -'sd38912;
    data[6239] = -'sd30719;
    data[6240] =  'sd10246;
    data[6241] =  'sd51230;
    data[6242] = -'sd71532;
    data[6243] = -'sd29978;
    data[6244] =  'sd13951;
    data[6245] =  'sd69755;
    data[6246] =  'sd21093;
    data[6247] = -'sd58376;
    data[6248] =  'sd35802;
    data[6249] =  'sd15169;
    data[6250] =  'sd75845;
    data[6251] =  'sd51543;
    data[6252] = -'sd69967;
    data[6253] = -'sd22153;
    data[6254] =  'sd53076;
    data[6255] = -'sd62302;
    data[6256] =  'sd16172;
    data[6257] =  'sd80860;
    data[6258] =  'sd76618;
    data[6259] =  'sd55408;
    data[6260] = -'sd50642;
    data[6261] =  'sd74472;
    data[6262] =  'sd44678;
    data[6263] =  'sd59549;
    data[6264] = -'sd29937;
    data[6265] =  'sd14156;
    data[6266] =  'sd70780;
    data[6267] =  'sd26218;
    data[6268] = -'sd32751;
    data[6269] =  'sd86;
    data[6270] =  'sd430;
    data[6271] =  'sd2150;
    data[6272] =  'sd10750;
    data[6273] =  'sd53750;
    data[6274] = -'sd58932;
    data[6275] =  'sd33022;
    data[6276] =  'sd1269;
    data[6277] =  'sd6345;
    data[6278] =  'sd31725;
    data[6279] = -'sd5216;
    data[6280] = -'sd26080;
    data[6281] =  'sd33441;
    data[6282] =  'sd3364;
    data[6283] =  'sd16820;
    data[6284] = -'sd79741;
    data[6285] = -'sd71023;
    data[6286] = -'sd27433;
    data[6287] =  'sd26676;
    data[6288] = -'sd30461;
    data[6289] =  'sd11536;
    data[6290] =  'sd57680;
    data[6291] = -'sd39282;
    data[6292] = -'sd32569;
    data[6293] =  'sd996;
    data[6294] =  'sd4980;
    data[6295] =  'sd24900;
    data[6296] = -'sd39341;
    data[6297] = -'sd32864;
    data[6298] = -'sd479;
    data[6299] = -'sd2395;
    data[6300] = -'sd11975;
    data[6301] = -'sd59875;
    data[6302] =  'sd28307;
    data[6303] = -'sd22306;
    data[6304] =  'sd52311;
    data[6305] = -'sd66127;
    data[6306] = -'sd2953;
    data[6307] = -'sd14765;
    data[6308] = -'sd73825;
    data[6309] = -'sd41443;
    data[6310] = -'sd43374;
    data[6311] = -'sd53029;
    data[6312] =  'sd62537;
    data[6313] = -'sd14997;
    data[6314] = -'sd74985;
    data[6315] = -'sd47243;
    data[6316] = -'sd72374;
    data[6317] = -'sd34188;
    data[6318] = -'sd7099;
    data[6319] = -'sd35495;
    data[6320] = -'sd13634;
    data[6321] = -'sd68170;
    data[6322] = -'sd13168;
    data[6323] = -'sd65840;
    data[6324] = -'sd1518;
    data[6325] = -'sd7590;
    data[6326] = -'sd37950;
    data[6327] = -'sd25909;
    data[6328] =  'sd34296;
    data[6329] =  'sd7639;
    data[6330] =  'sd38195;
    data[6331] =  'sd27134;
    data[6332] = -'sd28171;
    data[6333] =  'sd22986;
    data[6334] = -'sd48911;
    data[6335] = -'sd80714;
    data[6336] = -'sd75888;
    data[6337] = -'sd51758;
    data[6338] =  'sd68892;
    data[6339] =  'sd16778;
    data[6340] = -'sd79951;
    data[6341] = -'sd72073;
    data[6342] = -'sd32683;
    data[6343] =  'sd426;
    data[6344] =  'sd2130;
    data[6345] =  'sd10650;
    data[6346] =  'sd53250;
    data[6347] = -'sd61432;
    data[6348] =  'sd20522;
    data[6349] = -'sd61231;
    data[6350] =  'sd21527;
    data[6351] = -'sd56206;
    data[6352] =  'sd46652;
    data[6353] =  'sd69419;
    data[6354] =  'sd19413;
    data[6355] = -'sd66776;
    data[6356] = -'sd6198;
    data[6357] = -'sd30990;
    data[6358] =  'sd8891;
    data[6359] =  'sd44455;
    data[6360] =  'sd58434;
    data[6361] = -'sd35512;
    data[6362] = -'sd13719;
    data[6363] = -'sd68595;
    data[6364] = -'sd15293;
    data[6365] = -'sd76465;
    data[6366] = -'sd54643;
    data[6367] =  'sd54467;
    data[6368] = -'sd55347;
    data[6369] =  'sd50947;
    data[6370] = -'sd72947;
    data[6371] = -'sd37053;
    data[6372] = -'sd21424;
    data[6373] =  'sd56721;
    data[6374] = -'sd44077;
    data[6375] = -'sd56544;
    data[6376] =  'sd44962;
    data[6377] =  'sd60969;
    data[6378] = -'sd22837;
    data[6379] =  'sd49656;
    data[6380] = -'sd79402;
    data[6381] = -'sd69328;
    data[6382] = -'sd18958;
    data[6383] =  'sd69051;
    data[6384] =  'sd17573;
    data[6385] = -'sd75976;
    data[6386] = -'sd52198;
    data[6387] =  'sd66692;
    data[6388] =  'sd5778;
    data[6389] =  'sd28890;
    data[6390] = -'sd19391;
    data[6391] =  'sd66886;
    data[6392] =  'sd6748;
    data[6393] =  'sd33740;
    data[6394] =  'sd4859;
    data[6395] =  'sd24295;
    data[6396] = -'sd42366;
    data[6397] = -'sd47989;
    data[6398] = -'sd76104;
    data[6399] = -'sd52838;
    data[6400] =  'sd63492;
    data[6401] = -'sd10222;
    data[6402] = -'sd51110;
    data[6403] =  'sd72132;
    data[6404] =  'sd32978;
    data[6405] =  'sd1049;
    data[6406] =  'sd5245;
    data[6407] =  'sd26225;
    data[6408] = -'sd32716;
    data[6409] =  'sd261;
    data[6410] =  'sd1305;
    data[6411] =  'sd6525;
    data[6412] =  'sd32625;
    data[6413] = -'sd716;
    data[6414] = -'sd3580;
    data[6415] = -'sd17900;
    data[6416] =  'sd74341;
    data[6417] =  'sd44023;
    data[6418] =  'sd56274;
    data[6419] = -'sd46312;
    data[6420] = -'sd67719;
    data[6421] = -'sd10913;
    data[6422] = -'sd54565;
    data[6423] =  'sd54857;
    data[6424] = -'sd53397;
    data[6425] =  'sd60697;
    data[6426] = -'sd24197;
    data[6427] =  'sd42856;
    data[6428] =  'sd50439;
    data[6429] = -'sd75487;
    data[6430] = -'sd49753;
    data[6431] =  'sd78917;
    data[6432] =  'sd66903;
    data[6433] =  'sd6833;
    data[6434] =  'sd34165;
    data[6435] =  'sd6984;
    data[6436] =  'sd34920;
    data[6437] =  'sd10759;
    data[6438] =  'sd53795;
    data[6439] = -'sd58707;
    data[6440] =  'sd34147;
    data[6441] =  'sd6894;
    data[6442] =  'sd34470;
    data[6443] =  'sd8509;
    data[6444] =  'sd42545;
    data[6445] =  'sd48884;
    data[6446] =  'sd80579;
    data[6447] =  'sd75213;
    data[6448] =  'sd48383;
    data[6449] =  'sd78074;
    data[6450] =  'sd62688;
    data[6451] = -'sd14242;
    data[6452] = -'sd71210;
    data[6453] = -'sd28368;
    data[6454] =  'sd22001;
    data[6455] = -'sd53836;
    data[6456] =  'sd58502;
    data[6457] = -'sd35172;
    data[6458] = -'sd12019;
    data[6459] = -'sd60095;
    data[6460] =  'sd27207;
    data[6461] = -'sd27806;
    data[6462] =  'sd24811;
    data[6463] = -'sd39786;
    data[6464] = -'sd35089;
    data[6465] = -'sd11604;
    data[6466] = -'sd58020;
    data[6467] =  'sd37582;
    data[6468] =  'sd24069;
    data[6469] = -'sd43496;
    data[6470] = -'sd53639;
    data[6471] =  'sd59487;
    data[6472] = -'sd30247;
    data[6473] =  'sd12606;
    data[6474] =  'sd63030;
    data[6475] = -'sd12532;
    data[6476] = -'sd62660;
    data[6477] =  'sd14382;
    data[6478] =  'sd71910;
    data[6479] =  'sd31868;
    data[6480] = -'sd4501;
    data[6481] = -'sd22505;
    data[6482] =  'sd51316;
    data[6483] = -'sd71102;
    data[6484] = -'sd27828;
    data[6485] =  'sd24701;
    data[6486] = -'sd40336;
    data[6487] = -'sd37839;
    data[6488] = -'sd25354;
    data[6489] =  'sd37071;
    data[6490] =  'sd21514;
    data[6491] = -'sd56271;
    data[6492] =  'sd46327;
    data[6493] =  'sd67794;
    data[6494] =  'sd11288;
    data[6495] =  'sd56440;
    data[6496] = -'sd45482;
    data[6497] = -'sd63569;
    data[6498] =  'sd9837;
    data[6499] =  'sd49185;
    data[6500] = -'sd81757;
    data[6501] = -'sd81103;
    data[6502] = -'sd77833;
    data[6503] = -'sd61483;
    data[6504] =  'sd20267;
    data[6505] = -'sd62506;
    data[6506] =  'sd15152;
    data[6507] =  'sd75760;
    data[6508] =  'sd51118;
    data[6509] = -'sd72092;
    data[6510] = -'sd32778;
    data[6511] = -'sd49;
    data[6512] = -'sd245;
    data[6513] = -'sd1225;
    data[6514] = -'sd6125;
    data[6515] = -'sd30625;
    data[6516] =  'sd10716;
    data[6517] =  'sd53580;
    data[6518] = -'sd59782;
    data[6519] =  'sd28772;
    data[6520] = -'sd19981;
    data[6521] =  'sd63936;
    data[6522] = -'sd8002;
    data[6523] = -'sd40010;
    data[6524] = -'sd36209;
    data[6525] = -'sd17204;
    data[6526] =  'sd77821;
    data[6527] =  'sd61423;
    data[6528] = -'sd20567;
    data[6529] =  'sd61006;
    data[6530] = -'sd22652;
    data[6531] =  'sd50581;
    data[6532] = -'sd74777;
    data[6533] = -'sd46203;
    data[6534] = -'sd67174;
    data[6535] = -'sd8188;
    data[6536] = -'sd40940;
    data[6537] = -'sd40859;
    data[6538] = -'sd40454;
    data[6539] = -'sd38429;
    data[6540] = -'sd28304;
    data[6541] =  'sd22321;
    data[6542] = -'sd52236;
    data[6543] =  'sd66502;
    data[6544] =  'sd4828;
    data[6545] =  'sd24140;
    data[6546] = -'sd43141;
    data[6547] = -'sd51864;
    data[6548] =  'sd68362;
    data[6549] =  'sd14128;
    data[6550] =  'sd70640;
    data[6551] =  'sd25518;
    data[6552] = -'sd36251;
    data[6553] = -'sd17414;
    data[6554] =  'sd76771;
    data[6555] =  'sd56173;
    data[6556] = -'sd46817;
    data[6557] = -'sd70244;
    data[6558] = -'sd23538;
    data[6559] =  'sd46151;
    data[6560] =  'sd66914;
    data[6561] =  'sd6888;
    data[6562] =  'sd34440;
    data[6563] =  'sd8359;
    data[6564] =  'sd41795;
    data[6565] =  'sd45134;
    data[6566] =  'sd61829;
    data[6567] = -'sd18537;
    data[6568] =  'sd71156;
    data[6569] =  'sd28098;
    data[6570] = -'sd23351;
    data[6571] =  'sd47086;
    data[6572] =  'sd71589;
    data[6573] =  'sd30263;
    data[6574] = -'sd12526;
    data[6575] = -'sd62630;
    data[6576] =  'sd14532;
    data[6577] =  'sd72660;
    data[6578] =  'sd35618;
    data[6579] =  'sd14249;
    data[6580] =  'sd71245;
    data[6581] =  'sd28543;
    data[6582] = -'sd21126;
    data[6583] =  'sd58211;
    data[6584] = -'sd36627;
    data[6585] = -'sd19294;
    data[6586] =  'sd67371;
    data[6587] =  'sd9173;
    data[6588] =  'sd45865;
    data[6589] =  'sd65484;
    data[6590] = -'sd262;
    data[6591] = -'sd1310;
    data[6592] = -'sd6550;
    data[6593] = -'sd32750;
    data[6594] =  'sd91;
    data[6595] =  'sd455;
    data[6596] =  'sd2275;
    data[6597] =  'sd11375;
    data[6598] =  'sd56875;
    data[6599] = -'sd43307;
    data[6600] = -'sd52694;
    data[6601] =  'sd64212;
    data[6602] = -'sd6622;
    data[6603] = -'sd33110;
    data[6604] = -'sd1709;
    data[6605] = -'sd8545;
    data[6606] = -'sd42725;
    data[6607] = -'sd49784;
    data[6608] =  'sd78762;
    data[6609] =  'sd66128;
    data[6610] =  'sd2958;
    data[6611] =  'sd14790;
    data[6612] =  'sd73950;
    data[6613] =  'sd42068;
    data[6614] =  'sd46499;
    data[6615] =  'sd68654;
    data[6616] =  'sd15588;
    data[6617] =  'sd77940;
    data[6618] =  'sd62018;
    data[6619] = -'sd17592;
    data[6620] =  'sd75881;
    data[6621] =  'sd51723;
    data[6622] = -'sd69067;
    data[6623] = -'sd17653;
    data[6624] =  'sd75576;
    data[6625] =  'sd50198;
    data[6626] = -'sd76692;
    data[6627] = -'sd55778;
    data[6628] =  'sd48792;
    data[6629] =  'sd80119;
    data[6630] =  'sd72913;
    data[6631] =  'sd36883;
    data[6632] =  'sd20574;
    data[6633] = -'sd60971;
    data[6634] =  'sd22827;
    data[6635] = -'sd49706;
    data[6636] =  'sd79152;
    data[6637] =  'sd68078;
    data[6638] =  'sd12708;
    data[6639] =  'sd63540;
    data[6640] = -'sd9982;
    data[6641] = -'sd49910;
    data[6642] =  'sd78132;
    data[6643] =  'sd62978;
    data[6644] = -'sd12792;
    data[6645] = -'sd63960;
    data[6646] =  'sd7882;
    data[6647] =  'sd39410;
    data[6648] =  'sd33209;
    data[6649] =  'sd2204;
    data[6650] =  'sd11020;
    data[6651] =  'sd55100;
    data[6652] = -'sd52182;
    data[6653] =  'sd66772;
    data[6654] =  'sd6178;
    data[6655] =  'sd30890;
    data[6656] = -'sd9391;
    data[6657] = -'sd46955;
    data[6658] = -'sd70934;
    data[6659] = -'sd26988;
    data[6660] =  'sd28901;
    data[6661] = -'sd19336;
    data[6662] =  'sd67161;
    data[6663] =  'sd8123;
    data[6664] =  'sd40615;
    data[6665] =  'sd39234;
    data[6666] =  'sd32329;
    data[6667] = -'sd2196;
    data[6668] = -'sd10980;
    data[6669] = -'sd54900;
    data[6670] =  'sd53182;
    data[6671] = -'sd61772;
    data[6672] =  'sd18822;
    data[6673] = -'sd69731;
    data[6674] = -'sd20973;
    data[6675] =  'sd58976;
    data[6676] = -'sd32802;
    data[6677] = -'sd169;
    data[6678] = -'sd845;
    data[6679] = -'sd4225;
    data[6680] = -'sd21125;
    data[6681] =  'sd58216;
    data[6682] = -'sd36602;
    data[6683] = -'sd19169;
    data[6684] =  'sd67996;
    data[6685] =  'sd12298;
    data[6686] =  'sd61490;
    data[6687] = -'sd20232;
    data[6688] =  'sd62681;
    data[6689] = -'sd14277;
    data[6690] = -'sd71385;
    data[6691] = -'sd29243;
    data[6692] =  'sd17626;
    data[6693] = -'sd75711;
    data[6694] = -'sd50873;
    data[6695] =  'sd73317;
    data[6696] =  'sd38903;
    data[6697] =  'sd30674;
    data[6698] = -'sd10471;
    data[6699] = -'sd52355;
    data[6700] =  'sd65907;
    data[6701] =  'sd1853;
    data[6702] =  'sd9265;
    data[6703] =  'sd46325;
    data[6704] =  'sd67784;
    data[6705] =  'sd11238;
    data[6706] =  'sd56190;
    data[6707] = -'sd46732;
    data[6708] = -'sd69819;
    data[6709] = -'sd21413;
    data[6710] =  'sd56776;
    data[6711] = -'sd43802;
    data[6712] = -'sd55169;
    data[6713] =  'sd51837;
    data[6714] = -'sd68497;
    data[6715] = -'sd14803;
    data[6716] = -'sd74015;
    data[6717] = -'sd42393;
    data[6718] = -'sd48124;
    data[6719] = -'sd76779;
    data[6720] = -'sd56213;
    data[6721] =  'sd46617;
    data[6722] =  'sd69244;
    data[6723] =  'sd18538;
    data[6724] = -'sd71151;
    data[6725] = -'sd28073;
    data[6726] =  'sd23476;
    data[6727] = -'sd46461;
    data[6728] = -'sd68464;
    data[6729] = -'sd14638;
    data[6730] = -'sd73190;
    data[6731] = -'sd38268;
    data[6732] = -'sd27499;
    data[6733] =  'sd26346;
    data[6734] = -'sd32111;
    data[6735] =  'sd3286;
    data[6736] =  'sd16430;
    data[6737] = -'sd81691;
    data[6738] = -'sd80773;
    data[6739] = -'sd76183;
    data[6740] = -'sd53233;
    data[6741] =  'sd61517;
    data[6742] = -'sd20097;
    data[6743] =  'sd63356;
    data[6744] = -'sd10902;
    data[6745] = -'sd54510;
    data[6746] =  'sd55132;
    data[6747] = -'sd52022;
    data[6748] =  'sd67572;
    data[6749] =  'sd10178;
    data[6750] =  'sd50890;
    data[6751] = -'sd73232;
    data[6752] = -'sd38478;
    data[6753] = -'sd28549;
    data[6754] =  'sd21096;
    data[6755] = -'sd58361;
    data[6756] =  'sd35877;
    data[6757] =  'sd15544;
    data[6758] =  'sd77720;
    data[6759] =  'sd60918;
    data[6760] = -'sd23092;
    data[6761] =  'sd48381;
    data[6762] =  'sd78064;
    data[6763] =  'sd62638;
    data[6764] = -'sd14492;
    data[6765] = -'sd72460;
    data[6766] = -'sd34618;
    data[6767] = -'sd9249;
    data[6768] = -'sd46245;
    data[6769] = -'sd67384;
    data[6770] = -'sd9238;
    data[6771] = -'sd46190;
    data[6772] = -'sd67109;
    data[6773] = -'sd7863;
    data[6774] = -'sd39315;
    data[6775] = -'sd32734;
    data[6776] =  'sd171;
    data[6777] =  'sd855;
    data[6778] =  'sd4275;
    data[6779] =  'sd21375;
    data[6780] = -'sd56966;
    data[6781] =  'sd42852;
    data[6782] =  'sd50419;
    data[6783] = -'sd75587;
    data[6784] = -'sd50253;
    data[6785] =  'sd76417;
    data[6786] =  'sd54403;
    data[6787] = -'sd55667;
    data[6788] =  'sd49347;
    data[6789] = -'sd80947;
    data[6790] = -'sd77053;
    data[6791] = -'sd57583;
    data[6792] =  'sd39767;
    data[6793] =  'sd34994;
    data[6794] =  'sd11129;
    data[6795] =  'sd55645;
    data[6796] = -'sd49457;
    data[6797] =  'sd80397;
    data[6798] =  'sd74303;
    data[6799] =  'sd43833;
    data[6800] =  'sd55324;
    data[6801] = -'sd51062;
    data[6802] =  'sd72372;
    data[6803] =  'sd34178;
    data[6804] =  'sd7049;
    data[6805] =  'sd35245;
    data[6806] =  'sd12384;
    data[6807] =  'sd61920;
    data[6808] = -'sd18082;
    data[6809] =  'sd73431;
    data[6810] =  'sd39473;
    data[6811] =  'sd33524;
    data[6812] =  'sd3779;
    data[6813] =  'sd18895;
    data[6814] = -'sd69366;
    data[6815] = -'sd19148;
    data[6816] =  'sd68101;
    data[6817] =  'sd12823;
    data[6818] =  'sd64115;
    data[6819] = -'sd7107;
    data[6820] = -'sd35535;
    data[6821] = -'sd13834;
    data[6822] = -'sd69170;
    data[6823] = -'sd18168;
    data[6824] =  'sd73001;
    data[6825] =  'sd37323;
    data[6826] =  'sd22774;
    data[6827] = -'sd49971;
    data[6828] =  'sd77827;
    data[6829] =  'sd61453;
    data[6830] = -'sd20417;
    data[6831] =  'sd61756;
    data[6832] = -'sd18902;
    data[6833] =  'sd69331;
    data[6834] =  'sd18973;
    data[6835] = -'sd68976;
    data[6836] = -'sd17198;
    data[6837] =  'sd77851;
    data[6838] =  'sd61573;
    data[6839] = -'sd19817;
    data[6840] =  'sd64756;
    data[6841] = -'sd3902;
    data[6842] = -'sd19510;
    data[6843] =  'sd66291;
    data[6844] =  'sd3773;
    data[6845] =  'sd18865;
    data[6846] = -'sd69516;
    data[6847] = -'sd19898;
    data[6848] =  'sd64351;
    data[6849] = -'sd5927;
    data[6850] = -'sd29635;
    data[6851] =  'sd15666;
    data[6852] =  'sd78330;
    data[6853] =  'sd63968;
    data[6854] = -'sd7842;
    data[6855] = -'sd39210;
    data[6856] = -'sd32209;
    data[6857] =  'sd2796;
    data[6858] =  'sd13980;
    data[6859] =  'sd69900;
    data[6860] =  'sd21818;
    data[6861] = -'sd54751;
    data[6862] =  'sd53927;
    data[6863] = -'sd58047;
    data[6864] =  'sd37447;
    data[6865] =  'sd23394;
    data[6866] = -'sd46871;
    data[6867] = -'sd70514;
    data[6868] = -'sd24888;
    data[6869] =  'sd39401;
    data[6870] =  'sd33164;
    data[6871] =  'sd1979;
    data[6872] =  'sd9895;
    data[6873] =  'sd49475;
    data[6874] = -'sd80307;
    data[6875] = -'sd73853;
    data[6876] = -'sd41583;
    data[6877] = -'sd44074;
    data[6878] = -'sd56529;
    data[6879] =  'sd45037;
    data[6880] =  'sd61344;
    data[6881] = -'sd20962;
    data[6882] =  'sd59031;
    data[6883] = -'sd32527;
    data[6884] =  'sd1206;
    data[6885] =  'sd6030;
    data[6886] =  'sd30150;
    data[6887] = -'sd13091;
    data[6888] = -'sd65455;
    data[6889] =  'sd407;
    data[6890] =  'sd2035;
    data[6891] =  'sd10175;
    data[6892] =  'sd50875;
    data[6893] = -'sd73307;
    data[6894] = -'sd38853;
    data[6895] = -'sd30424;
    data[6896] =  'sd11721;
    data[6897] =  'sd58605;
    data[6898] = -'sd34657;
    data[6899] = -'sd9444;
    data[6900] = -'sd47220;
    data[6901] = -'sd72259;
    data[6902] = -'sd33613;
    data[6903] = -'sd4224;
    data[6904] = -'sd21120;
    data[6905] =  'sd58241;
    data[6906] = -'sd36477;
    data[6907] = -'sd18544;
    data[6908] =  'sd71121;
    data[6909] =  'sd27923;
    data[6910] = -'sd24226;
    data[6911] =  'sd42711;
    data[6912] =  'sd49714;
    data[6913] = -'sd79112;
    data[6914] = -'sd67878;
    data[6915] = -'sd11708;
    data[6916] = -'sd58540;
    data[6917] =  'sd34982;
    data[6918] =  'sd11069;
    data[6919] =  'sd55345;
    data[6920] = -'sd50957;
    data[6921] =  'sd72897;
    data[6922] =  'sd36803;
    data[6923] =  'sd20174;
    data[6924] = -'sd62971;
    data[6925] =  'sd12827;
    data[6926] =  'sd64135;
    data[6927] = -'sd7007;
    data[6928] = -'sd35035;
    data[6929] = -'sd11334;
    data[6930] = -'sd56670;
    data[6931] =  'sd44332;
    data[6932] =  'sd57819;
    data[6933] = -'sd38587;
    data[6934] = -'sd29094;
    data[6935] =  'sd18371;
    data[6936] = -'sd71986;
    data[6937] = -'sd32248;
    data[6938] =  'sd2601;
    data[6939] =  'sd13005;
    data[6940] =  'sd65025;
    data[6941] = -'sd2557;
    data[6942] = -'sd12785;
    data[6943] = -'sd63925;
    data[6944] =  'sd8057;
    data[6945] =  'sd40285;
    data[6946] =  'sd37584;
    data[6947] =  'sd24079;
    data[6948] = -'sd43446;
    data[6949] = -'sd53389;
    data[6950] =  'sd60737;
    data[6951] = -'sd23997;
    data[6952] =  'sd43856;
    data[6953] =  'sd55439;
    data[6954] = -'sd50487;
    data[6955] =  'sd75247;
    data[6956] =  'sd48553;
    data[6957] =  'sd78924;
    data[6958] =  'sd66938;
    data[6959] =  'sd7008;
    data[6960] =  'sd35040;
    data[6961] =  'sd11359;
    data[6962] =  'sd56795;
    data[6963] = -'sd43707;
    data[6964] = -'sd54694;
    data[6965] =  'sd54212;
    data[6966] = -'sd56622;
    data[6967] =  'sd44572;
    data[6968] =  'sd59019;
    data[6969] = -'sd32587;
    data[6970] =  'sd906;
    data[6971] =  'sd4530;
    data[6972] =  'sd22650;
    data[6973] = -'sd50591;
    data[6974] =  'sd74727;
    data[6975] =  'sd45953;
    data[6976] =  'sd65924;
    data[6977] =  'sd1938;
    data[6978] =  'sd9690;
    data[6979] =  'sd48450;
    data[6980] =  'sd78409;
    data[6981] =  'sd64363;
    data[6982] = -'sd5867;
    data[6983] = -'sd29335;
    data[6984] =  'sd17166;
    data[6985] = -'sd78011;
    data[6986] = -'sd62373;
    data[6987] =  'sd15817;
    data[6988] =  'sd79085;
    data[6989] =  'sd67743;
    data[6990] =  'sd11033;
    data[6991] =  'sd55165;
    data[6992] = -'sd51857;
    data[6993] =  'sd68397;
    data[6994] =  'sd14303;
    data[6995] =  'sd71515;
    data[6996] =  'sd29893;
    data[6997] = -'sd14376;
    data[6998] = -'sd71880;
    data[6999] = -'sd31718;
    data[7000] =  'sd5251;
    data[7001] =  'sd26255;
    data[7002] = -'sd32566;
    data[7003] =  'sd1011;
    data[7004] =  'sd5055;
    data[7005] =  'sd25275;
    data[7006] = -'sd37466;
    data[7007] = -'sd23489;
    data[7008] =  'sd46396;
    data[7009] =  'sd68139;
    data[7010] =  'sd13013;
    data[7011] =  'sd65065;
    data[7012] = -'sd2357;
    data[7013] = -'sd11785;
    data[7014] = -'sd58925;
    data[7015] =  'sd33057;
    data[7016] =  'sd1444;
    data[7017] =  'sd7220;
    data[7018] =  'sd36100;
    data[7019] =  'sd16659;
    data[7020] = -'sd80546;
    data[7021] = -'sd75048;
    data[7022] = -'sd47558;
    data[7023] = -'sd73949;
    data[7024] = -'sd42063;
    data[7025] = -'sd46474;
    data[7026] = -'sd68529;
    data[7027] = -'sd14963;
    data[7028] = -'sd74815;
    data[7029] = -'sd46393;
    data[7030] = -'sd68124;
    data[7031] = -'sd12938;
    data[7032] = -'sd64690;
    data[7033] =  'sd4232;
    data[7034] =  'sd21160;
    data[7035] = -'sd58041;
    data[7036] =  'sd37477;
    data[7037] =  'sd23544;
    data[7038] = -'sd46121;
    data[7039] = -'sd66764;
    data[7040] = -'sd6138;
    data[7041] = -'sd30690;
    data[7042] =  'sd10391;
    data[7043] =  'sd51955;
    data[7044] = -'sd67907;
    data[7045] = -'sd11853;
    data[7046] = -'sd59265;
    data[7047] =  'sd31357;
    data[7048] = -'sd7056;
    data[7049] = -'sd35280;
    data[7050] = -'sd12559;
    data[7051] = -'sd62795;
    data[7052] =  'sd13707;
    data[7053] =  'sd68535;
    data[7054] =  'sd14993;
    data[7055] =  'sd74965;
    data[7056] =  'sd47143;
    data[7057] =  'sd71874;
    data[7058] =  'sd31688;
    data[7059] = -'sd5401;
    data[7060] = -'sd27005;
    data[7061] =  'sd28816;
    data[7062] = -'sd19761;
    data[7063] =  'sd65036;
    data[7064] = -'sd2502;
    data[7065] = -'sd12510;
    data[7066] = -'sd62550;
    data[7067] =  'sd14932;
    data[7068] =  'sd74660;
    data[7069] =  'sd45618;
    data[7070] =  'sd64249;
    data[7071] = -'sd6437;
    data[7072] = -'sd32185;
    data[7073] =  'sd2916;
    data[7074] =  'sd14580;
    data[7075] =  'sd72900;
    data[7076] =  'sd36818;
    data[7077] =  'sd20249;
    data[7078] = -'sd62596;
    data[7079] =  'sd14702;
    data[7080] =  'sd73510;
    data[7081] =  'sd39868;
    data[7082] =  'sd35499;
    data[7083] =  'sd13654;
    data[7084] =  'sd68270;
    data[7085] =  'sd13668;
    data[7086] =  'sd68340;
    data[7087] =  'sd14018;
    data[7088] =  'sd70090;
    data[7089] =  'sd22768;
    data[7090] = -'sd50001;
    data[7091] =  'sd77677;
    data[7092] =  'sd60703;
    data[7093] = -'sd24167;
    data[7094] =  'sd43006;
    data[7095] =  'sd51189;
    data[7096] = -'sd71737;
    data[7097] = -'sd31003;
    data[7098] =  'sd8826;
    data[7099] =  'sd44130;
    data[7100] =  'sd56809;
    data[7101] = -'sd43637;
    data[7102] = -'sd54344;
    data[7103] =  'sd55962;
    data[7104] = -'sd47872;
    data[7105] = -'sd75519;
    data[7106] = -'sd49913;
    data[7107] =  'sd78117;
    data[7108] =  'sd62903;
    data[7109] = -'sd13167;
    data[7110] = -'sd65835;
    data[7111] = -'sd1493;
    data[7112] = -'sd7465;
    data[7113] = -'sd37325;
    data[7114] = -'sd22784;
    data[7115] =  'sd49921;
    data[7116] = -'sd78077;
    data[7117] = -'sd62703;
    data[7118] =  'sd14167;
    data[7119] =  'sd70835;
    data[7120] =  'sd26493;
    data[7121] = -'sd31376;
    data[7122] =  'sd6961;
    data[7123] =  'sd34805;
    data[7124] =  'sd10184;
    data[7125] =  'sd50920;
    data[7126] = -'sd73082;
    data[7127] = -'sd37728;
    data[7128] = -'sd24799;
    data[7129] =  'sd39846;
    data[7130] =  'sd35389;
    data[7131] =  'sd13104;
    data[7132] =  'sd65520;
    data[7133] = -'sd82;
    data[7134] = -'sd410;
    data[7135] = -'sd2050;
    data[7136] = -'sd10250;
    data[7137] = -'sd51250;
    data[7138] =  'sd71432;
    data[7139] =  'sd29478;
    data[7140] = -'sd16451;
    data[7141] =  'sd81586;
    data[7142] =  'sd80248;
    data[7143] =  'sd73558;
    data[7144] =  'sd40108;
    data[7145] =  'sd36699;
    data[7146] =  'sd19654;
    data[7147] = -'sd65571;
    data[7148] = -'sd173;
    data[7149] = -'sd865;
    data[7150] = -'sd4325;
    data[7151] = -'sd21625;
    data[7152] =  'sd55716;
    data[7153] = -'sd49102;
    data[7154] = -'sd81669;
    data[7155] = -'sd80663;
    data[7156] = -'sd75633;
    data[7157] = -'sd50483;
    data[7158] =  'sd75267;
    data[7159] =  'sd48653;
    data[7160] =  'sd79424;
    data[7161] =  'sd69438;
    data[7162] =  'sd19508;
    data[7163] = -'sd66301;
    data[7164] = -'sd3823;
    data[7165] = -'sd19115;
    data[7166] =  'sd68266;
    data[7167] =  'sd13648;
    data[7168] =  'sd68240;
    data[7169] =  'sd13518;
    data[7170] =  'sd67590;
    data[7171] =  'sd10268;
    data[7172] =  'sd51340;
    data[7173] = -'sd70982;
    data[7174] = -'sd27228;
    data[7175] =  'sd27701;
    data[7176] = -'sd25336;
    data[7177] =  'sd37161;
    data[7178] =  'sd21964;
    data[7179] = -'sd54021;
    data[7180] =  'sd57577;
    data[7181] = -'sd39797;
    data[7182] = -'sd35144;
    data[7183] = -'sd11879;
    data[7184] = -'sd59395;
    data[7185] =  'sd30707;
    data[7186] = -'sd10306;
    data[7187] = -'sd51530;
    data[7188] =  'sd70032;
    data[7189] =  'sd22478;
    data[7190] = -'sd51451;
    data[7191] =  'sd70427;
    data[7192] =  'sd24453;
    data[7193] = -'sd41576;
    data[7194] = -'sd44039;
    data[7195] = -'sd56354;
    data[7196] =  'sd45912;
    data[7197] =  'sd65719;
    data[7198] =  'sd913;
    data[7199] =  'sd4565;
    data[7200] =  'sd22825;
    data[7201] = -'sd49716;
    data[7202] =  'sd79102;
    data[7203] =  'sd67828;
    data[7204] =  'sd11458;
    data[7205] =  'sd57290;
    data[7206] = -'sd41232;
    data[7207] = -'sd42319;
    data[7208] = -'sd47754;
    data[7209] = -'sd74929;
    data[7210] = -'sd46963;
    data[7211] = -'sd70974;
    data[7212] = -'sd27188;
    data[7213] =  'sd27901;
    data[7214] = -'sd24336;
    data[7215] =  'sd42161;
    data[7216] =  'sd46964;
    data[7217] =  'sd70979;
    data[7218] =  'sd27213;
    data[7219] = -'sd27776;
    data[7220] =  'sd24961;
    data[7221] = -'sd39036;
    data[7222] = -'sd31339;
    data[7223] =  'sd7146;
    data[7224] =  'sd35730;
    data[7225] =  'sd14809;
    data[7226] =  'sd74045;
    data[7227] =  'sd42543;
    data[7228] =  'sd48874;
    data[7229] =  'sd80529;
    data[7230] =  'sd74963;
    data[7231] =  'sd47133;
    data[7232] =  'sd71824;
    data[7233] =  'sd31438;
    data[7234] = -'sd6651;
    data[7235] = -'sd33255;
    data[7236] = -'sd2434;
    data[7237] = -'sd12170;
    data[7238] = -'sd60850;
    data[7239] =  'sd23432;
    data[7240] = -'sd46681;
    data[7241] = -'sd69564;
    data[7242] = -'sd20138;
    data[7243] =  'sd63151;
    data[7244] = -'sd11927;
    data[7245] = -'sd59635;
    data[7246] =  'sd29507;
    data[7247] = -'sd16306;
    data[7248] = -'sd81530;
    data[7249] = -'sd79968;
    data[7250] = -'sd72158;
    data[7251] = -'sd33108;
    data[7252] = -'sd1699;
    data[7253] = -'sd8495;
    data[7254] = -'sd42475;
    data[7255] = -'sd48534;
    data[7256] = -'sd78829;
    data[7257] = -'sd66463;
    data[7258] = -'sd4633;
    data[7259] = -'sd23165;
    data[7260] =  'sd48016;
    data[7261] =  'sd76239;
    data[7262] =  'sd53513;
    data[7263] = -'sd60117;
    data[7264] =  'sd27097;
    data[7265] = -'sd28356;
    data[7266] =  'sd22061;
    data[7267] = -'sd53536;
    data[7268] =  'sd60002;
    data[7269] = -'sd27672;
    data[7270] =  'sd25481;
    data[7271] = -'sd36436;
    data[7272] = -'sd18339;
    data[7273] =  'sd72146;
    data[7274] =  'sd33048;
    data[7275] =  'sd1399;
    data[7276] =  'sd6995;
    data[7277] =  'sd34975;
    data[7278] =  'sd11034;
    data[7279] =  'sd55170;
    data[7280] = -'sd51832;
    data[7281] =  'sd68522;
    data[7282] =  'sd14928;
    data[7283] =  'sd74640;
    data[7284] =  'sd45518;
    data[7285] =  'sd63749;
    data[7286] = -'sd8937;
    data[7287] = -'sd44685;
    data[7288] = -'sd59584;
    data[7289] =  'sd29762;
    data[7290] = -'sd15031;
    data[7291] = -'sd75155;
    data[7292] = -'sd48093;
    data[7293] = -'sd76624;
    data[7294] = -'sd55438;
    data[7295] =  'sd50492;
    data[7296] = -'sd75222;
    data[7297] = -'sd48428;
    data[7298] = -'sd78299;
    data[7299] = -'sd63813;
    data[7300] =  'sd8617;
    data[7301] =  'sd43085;
    data[7302] =  'sd51584;
    data[7303] = -'sd69762;
    data[7304] = -'sd21128;
    data[7305] =  'sd58201;
    data[7306] = -'sd36677;
    data[7307] = -'sd19544;
    data[7308] =  'sd66121;
    data[7309] =  'sd2923;
    data[7310] =  'sd14615;
    data[7311] =  'sd73075;
    data[7312] =  'sd37693;
    data[7313] =  'sd24624;
    data[7314] = -'sd40721;
    data[7315] = -'sd39764;
    data[7316] = -'sd34979;
    data[7317] = -'sd11054;
    data[7318] = -'sd55270;
    data[7319] =  'sd51332;
    data[7320] = -'sd71022;
    data[7321] = -'sd27428;
    data[7322] =  'sd26701;
    data[7323] = -'sd30336;
    data[7324] =  'sd12161;
    data[7325] =  'sd60805;
    data[7326] = -'sd23657;
    data[7327] =  'sd45556;
    data[7328] =  'sd63939;
    data[7329] = -'sd7987;
    data[7330] = -'sd39935;
    data[7331] = -'sd35834;
    data[7332] = -'sd15329;
    data[7333] = -'sd76645;
    data[7334] = -'sd55543;
    data[7335] =  'sd49967;
    data[7336] = -'sd77847;
    data[7337] = -'sd61553;
    data[7338] =  'sd19917;
    data[7339] = -'sd64256;
    data[7340] =  'sd6402;
    data[7341] =  'sd32010;
    data[7342] = -'sd3791;
    data[7343] = -'sd18955;
    data[7344] =  'sd69066;
    data[7345] =  'sd17648;
    data[7346] = -'sd75601;
    data[7347] = -'sd50323;
    data[7348] =  'sd76067;
    data[7349] =  'sd52653;
    data[7350] = -'sd64417;
    data[7351] =  'sd5597;
    data[7352] =  'sd27985;
    data[7353] = -'sd23916;
    data[7354] =  'sd44261;
    data[7355] =  'sd57464;
    data[7356] = -'sd40362;
    data[7357] = -'sd37969;
    data[7358] = -'sd26004;
    data[7359] =  'sd33821;
    data[7360] =  'sd5264;
    data[7361] =  'sd26320;
    data[7362] = -'sd32241;
    data[7363] =  'sd2636;
    data[7364] =  'sd13180;
    data[7365] =  'sd65900;
    data[7366] =  'sd1818;
    data[7367] =  'sd9090;
    data[7368] =  'sd45450;
    data[7369] =  'sd63409;
    data[7370] = -'sd10637;
    data[7371] = -'sd53185;
    data[7372] =  'sd61757;
    data[7373] = -'sd18897;
    data[7374] =  'sd69356;
    data[7375] =  'sd19098;
    data[7376] = -'sd68351;
    data[7377] = -'sd14073;
    data[7378] = -'sd70365;
    data[7379] = -'sd24143;
    data[7380] =  'sd43126;
    data[7381] =  'sd51789;
    data[7382] = -'sd68737;
    data[7383] = -'sd16003;
    data[7384] = -'sd80015;
    data[7385] = -'sd72393;
    data[7386] = -'sd34283;
    data[7387] = -'sd7574;
    data[7388] = -'sd37870;
    data[7389] = -'sd25509;
    data[7390] =  'sd36296;
    data[7391] =  'sd17639;
    data[7392] = -'sd75646;
    data[7393] = -'sd50548;
    data[7394] =  'sd74942;
    data[7395] =  'sd47028;
    data[7396] =  'sd71299;
    data[7397] =  'sd28813;
    data[7398] = -'sd19776;
    data[7399] =  'sd64961;
    data[7400] = -'sd2877;
    data[7401] = -'sd14385;
    data[7402] = -'sd71925;
    data[7403] = -'sd31943;
    data[7404] =  'sd4126;
    data[7405] =  'sd20630;
    data[7406] = -'sd60691;
    data[7407] =  'sd24227;
    data[7408] = -'sd42706;
    data[7409] = -'sd49689;
    data[7410] =  'sd79237;
    data[7411] =  'sd68503;
    data[7412] =  'sd14833;
    data[7413] =  'sd74165;
    data[7414] =  'sd43143;
    data[7415] =  'sd51874;
    data[7416] = -'sd68312;
    data[7417] = -'sd13878;
    data[7418] = -'sd69390;
    data[7419] = -'sd19268;
    data[7420] =  'sd67501;
    data[7421] =  'sd9823;
    data[7422] =  'sd49115;
    data[7423] =  'sd81734;
    data[7424] =  'sd80988;
    data[7425] =  'sd77258;
    data[7426] =  'sd58608;
    data[7427] = -'sd34642;
    data[7428] = -'sd9369;
    data[7429] = -'sd46845;
    data[7430] = -'sd70384;
    data[7431] = -'sd24238;
    data[7432] =  'sd42651;
    data[7433] =  'sd49414;
    data[7434] = -'sd80612;
    data[7435] = -'sd75378;
    data[7436] = -'sd49208;
    data[7437] =  'sd81642;
    data[7438] =  'sd80528;
    data[7439] =  'sd74958;
    data[7440] =  'sd47108;
    data[7441] =  'sd71699;
    data[7442] =  'sd30813;
    data[7443] = -'sd9776;
    data[7444] = -'sd48880;
    data[7445] = -'sd80559;
    data[7446] = -'sd75113;
    data[7447] = -'sd47883;
    data[7448] = -'sd75574;
    data[7449] = -'sd50188;
    data[7450] =  'sd76742;
    data[7451] =  'sd56028;
    data[7452] = -'sd47542;
    data[7453] = -'sd73869;
    data[7454] = -'sd41663;
    data[7455] = -'sd44474;
    data[7456] = -'sd58529;
    data[7457] =  'sd35037;
    data[7458] =  'sd11344;
    data[7459] =  'sd56720;
    data[7460] = -'sd44082;
    data[7461] = -'sd56569;
    data[7462] =  'sd44837;
    data[7463] =  'sd60344;
    data[7464] = -'sd25962;
    data[7465] =  'sd34031;
    data[7466] =  'sd6314;
    data[7467] =  'sd31570;
    data[7468] = -'sd5991;
    data[7469] = -'sd29955;
    data[7470] =  'sd14066;
    data[7471] =  'sd70330;
    data[7472] =  'sd23968;
    data[7473] = -'sd44001;
    data[7474] = -'sd56164;
    data[7475] =  'sd46862;
    data[7476] =  'sd70469;
    data[7477] =  'sd24663;
    data[7478] = -'sd40526;
    data[7479] = -'sd38789;
    data[7480] = -'sd30104;
    data[7481] =  'sd13321;
    data[7482] =  'sd66605;
    data[7483] =  'sd5343;
    data[7484] =  'sd26715;
    data[7485] = -'sd30266;
    data[7486] =  'sd12511;
    data[7487] =  'sd62555;
    data[7488] = -'sd14907;
    data[7489] = -'sd74535;
    data[7490] = -'sd44993;
    data[7491] = -'sd61124;
    data[7492] =  'sd22062;
    data[7493] = -'sd53531;
    data[7494] =  'sd60027;
    data[7495] = -'sd27547;
    data[7496] =  'sd26106;
    data[7497] = -'sd33311;
    data[7498] = -'sd2714;
    data[7499] = -'sd13570;
    data[7500] = -'sd67850;
    data[7501] = -'sd11568;
    data[7502] = -'sd57840;
    data[7503] =  'sd38482;
    data[7504] =  'sd28569;
    data[7505] = -'sd20996;
    data[7506] =  'sd58861;
    data[7507] = -'sd33377;
    data[7508] = -'sd3044;
    data[7509] = -'sd15220;
    data[7510] = -'sd76100;
    data[7511] = -'sd52818;
    data[7512] =  'sd63592;
    data[7513] = -'sd9722;
    data[7514] = -'sd48610;
    data[7515] = -'sd79209;
    data[7516] = -'sd68363;
    data[7517] = -'sd14133;
    data[7518] = -'sd70665;
    data[7519] = -'sd25643;
    data[7520] =  'sd35626;
    data[7521] =  'sd14289;
    data[7522] =  'sd71445;
    data[7523] =  'sd29543;
    data[7524] = -'sd16126;
    data[7525] = -'sd80630;
    data[7526] = -'sd75468;
    data[7527] = -'sd49658;
    data[7528] =  'sd79392;
    data[7529] =  'sd69278;
    data[7530] =  'sd18708;
    data[7531] = -'sd70301;
    data[7532] = -'sd23823;
    data[7533] =  'sd44726;
    data[7534] =  'sd59789;
    data[7535] = -'sd28737;
    data[7536] =  'sd20156;
    data[7537] = -'sd63061;
    data[7538] =  'sd12377;
    data[7539] =  'sd61885;
    data[7540] = -'sd18257;
    data[7541] =  'sd72556;
    data[7542] =  'sd35098;
    data[7543] =  'sd11649;
    data[7544] =  'sd58245;
    data[7545] = -'sd36457;
    data[7546] = -'sd18444;
    data[7547] =  'sd71621;
    data[7548] =  'sd30423;
    data[7549] = -'sd11726;
    data[7550] = -'sd58630;
    data[7551] =  'sd34532;
    data[7552] =  'sd8819;
    data[7553] =  'sd44095;
    data[7554] =  'sd56634;
    data[7555] = -'sd44512;
    data[7556] = -'sd58719;
    data[7557] =  'sd34087;
    data[7558] =  'sd6594;
    data[7559] =  'sd32970;
    data[7560] =  'sd1009;
    data[7561] =  'sd5045;
    data[7562] =  'sd25225;
    data[7563] = -'sd37716;
    data[7564] = -'sd24739;
    data[7565] =  'sd40146;
    data[7566] =  'sd36889;
    data[7567] =  'sd20604;
    data[7568] = -'sd60821;
    data[7569] =  'sd23577;
    data[7570] = -'sd45956;
    data[7571] = -'sd65939;
    data[7572] = -'sd2013;
    data[7573] = -'sd10065;
    data[7574] = -'sd50325;
    data[7575] =  'sd76057;
    data[7576] =  'sd52603;
    data[7577] = -'sd64667;
    data[7578] =  'sd4347;
    data[7579] =  'sd21735;
    data[7580] = -'sd55166;
    data[7581] =  'sd51852;
    data[7582] = -'sd68422;
    data[7583] = -'sd14428;
    data[7584] = -'sd72140;
    data[7585] = -'sd33018;
    data[7586] = -'sd1249;
    data[7587] = -'sd6245;
    data[7588] = -'sd31225;
    data[7589] =  'sd7716;
    data[7590] =  'sd38580;
    data[7591] =  'sd29059;
    data[7592] = -'sd18546;
    data[7593] =  'sd71111;
    data[7594] =  'sd27873;
    data[7595] = -'sd24476;
    data[7596] =  'sd41461;
    data[7597] =  'sd43464;
    data[7598] =  'sd53479;
    data[7599] = -'sd60287;
    data[7600] =  'sd26247;
    data[7601] = -'sd32606;
    data[7602] =  'sd811;
    data[7603] =  'sd4055;
    data[7604] =  'sd20275;
    data[7605] = -'sd62466;
    data[7606] =  'sd15352;
    data[7607] =  'sd76760;
    data[7608] =  'sd56118;
    data[7609] = -'sd47092;
    data[7610] = -'sd71619;
    data[7611] = -'sd30413;
    data[7612] =  'sd11776;
    data[7613] =  'sd58880;
    data[7614] = -'sd33282;
    data[7615] = -'sd2569;
    data[7616] = -'sd12845;
    data[7617] = -'sd64225;
    data[7618] =  'sd6557;
    data[7619] =  'sd32785;
    data[7620] =  'sd84;
    data[7621] =  'sd420;
    data[7622] =  'sd2100;
    data[7623] =  'sd10500;
    data[7624] =  'sd52500;
    data[7625] = -'sd65182;
    data[7626] =  'sd1772;
    data[7627] =  'sd8860;
    data[7628] =  'sd44300;
    data[7629] =  'sd57659;
    data[7630] = -'sd39387;
    data[7631] = -'sd33094;
    data[7632] = -'sd1629;
    data[7633] = -'sd8145;
    data[7634] = -'sd40725;
    data[7635] = -'sd39784;
    data[7636] = -'sd35079;
    data[7637] = -'sd11554;
    data[7638] = -'sd57770;
    data[7639] =  'sd38832;
    data[7640] =  'sd30319;
    data[7641] = -'sd12246;
    data[7642] = -'sd61230;
    data[7643] =  'sd21532;
    data[7644] = -'sd56181;
    data[7645] =  'sd46777;
    data[7646] =  'sd70044;
    data[7647] =  'sd22538;
    data[7648] = -'sd51151;
    data[7649] =  'sd71927;
    data[7650] =  'sd31953;
    data[7651] = -'sd4076;
    data[7652] = -'sd20380;
    data[7653] =  'sd61941;
    data[7654] = -'sd17977;
    data[7655] =  'sd73956;
    data[7656] =  'sd42098;
    data[7657] =  'sd46649;
    data[7658] =  'sd69404;
    data[7659] =  'sd19338;
    data[7660] = -'sd67151;
    data[7661] = -'sd8073;
    data[7662] = -'sd40365;
    data[7663] = -'sd37984;
    data[7664] = -'sd26079;
    data[7665] =  'sd33446;
    data[7666] =  'sd3389;
    data[7667] =  'sd16945;
    data[7668] = -'sd79116;
    data[7669] = -'sd67898;
    data[7670] = -'sd11808;
    data[7671] = -'sd59040;
    data[7672] =  'sd32482;
    data[7673] = -'sd1431;
    data[7674] = -'sd7155;
    data[7675] = -'sd35775;
    data[7676] = -'sd15034;
    data[7677] = -'sd75170;
    data[7678] = -'sd48168;
    data[7679] = -'sd76999;
    data[7680] = -'sd57313;
    data[7681] =  'sd41117;
    data[7682] =  'sd41744;
    data[7683] =  'sd44879;
    data[7684] =  'sd60554;
    data[7685] = -'sd24912;
    data[7686] =  'sd39281;
    data[7687] =  'sd32564;
    data[7688] = -'sd1021;
    data[7689] = -'sd5105;
    data[7690] = -'sd25525;
    data[7691] =  'sd36216;
    data[7692] =  'sd17239;
    data[7693] = -'sd77646;
    data[7694] = -'sd60548;
    data[7695] =  'sd24942;
    data[7696] = -'sd39131;
    data[7697] = -'sd31814;
    data[7698] =  'sd4771;
    data[7699] =  'sd23855;
    data[7700] = -'sd44566;
    data[7701] = -'sd58989;
    data[7702] =  'sd32737;
    data[7703] = -'sd156;
    data[7704] = -'sd780;
    data[7705] = -'sd3900;
    data[7706] = -'sd19500;
    data[7707] =  'sd66341;
    data[7708] =  'sd4023;
    data[7709] =  'sd20115;
    data[7710] = -'sd63266;
    data[7711] =  'sd11352;
    data[7712] =  'sd56760;
    data[7713] = -'sd43882;
    data[7714] = -'sd55569;
    data[7715] =  'sd49837;
    data[7716] = -'sd78497;
    data[7717] = -'sd64803;
    data[7718] =  'sd3667;
    data[7719] =  'sd18335;
    data[7720] = -'sd72166;
    data[7721] = -'sd33148;
    data[7722] = -'sd1899;
    data[7723] = -'sd9495;
    data[7724] = -'sd47475;
    data[7725] = -'sd73534;
    data[7726] = -'sd39988;
    data[7727] = -'sd36099;
    data[7728] = -'sd16654;
    data[7729] =  'sd80571;
    data[7730] =  'sd75173;
    data[7731] =  'sd48183;
    data[7732] =  'sd77074;
    data[7733] =  'sd57688;
    data[7734] = -'sd39242;
    data[7735] = -'sd32369;
    data[7736] =  'sd1996;
    data[7737] =  'sd9980;
    data[7738] =  'sd49900;
    data[7739] = -'sd78182;
    data[7740] = -'sd63228;
    data[7741] =  'sd11542;
    data[7742] =  'sd57710;
    data[7743] = -'sd39132;
    data[7744] = -'sd31819;
    data[7745] =  'sd4746;
    data[7746] =  'sd23730;
    data[7747] = -'sd45191;
    data[7748] = -'sd62114;
    data[7749] =  'sd17112;
    data[7750] = -'sd78281;
    data[7751] = -'sd63723;
    data[7752] =  'sd9067;
    data[7753] =  'sd45335;
    data[7754] =  'sd62834;
    data[7755] = -'sd13512;
    data[7756] = -'sd67560;
    data[7757] = -'sd10118;
    data[7758] = -'sd50590;
    data[7759] =  'sd74732;
    data[7760] =  'sd45978;
    data[7761] =  'sd66049;
    data[7762] =  'sd2563;
    data[7763] =  'sd12815;
    data[7764] =  'sd64075;
    data[7765] = -'sd7307;
    data[7766] = -'sd36535;
    data[7767] = -'sd18834;
    data[7768] =  'sd69671;
    data[7769] =  'sd20673;
    data[7770] = -'sd60476;
    data[7771] =  'sd25302;
    data[7772] = -'sd37331;
    data[7773] = -'sd22814;
    data[7774] =  'sd49771;
    data[7775] = -'sd78827;
    data[7776] = -'sd66453;
    data[7777] = -'sd4583;
    data[7778] = -'sd22915;
    data[7779] =  'sd49266;
    data[7780] = -'sd81352;
    data[7781] = -'sd79078;
    data[7782] = -'sd67708;
    data[7783] = -'sd10858;
    data[7784] = -'sd54290;
    data[7785] =  'sd56232;
    data[7786] = -'sd46522;
    data[7787] = -'sd68769;
    data[7788] = -'sd16163;
    data[7789] = -'sd80815;
    data[7790] = -'sd76393;
    data[7791] = -'sd54283;
    data[7792] =  'sd56267;
    data[7793] = -'sd46347;
    data[7794] = -'sd67894;
    data[7795] = -'sd11788;
    data[7796] = -'sd58940;
    data[7797] =  'sd32982;
    data[7798] =  'sd1069;
    data[7799] =  'sd5345;
    data[7800] =  'sd26725;
    data[7801] = -'sd30216;
    data[7802] =  'sd12761;
    data[7803] =  'sd63805;
    data[7804] = -'sd8657;
    data[7805] = -'sd43285;
    data[7806] = -'sd52584;
    data[7807] =  'sd64762;
    data[7808] = -'sd3872;
    data[7809] = -'sd19360;
    data[7810] =  'sd67041;
    data[7811] =  'sd7523;
    data[7812] =  'sd37615;
    data[7813] =  'sd24234;
    data[7814] = -'sd42671;
    data[7815] = -'sd49514;
    data[7816] =  'sd80112;
    data[7817] =  'sd72878;
    data[7818] =  'sd36708;
    data[7819] =  'sd19699;
    data[7820] = -'sd65346;
    data[7821] =  'sd952;
    data[7822] =  'sd4760;
    data[7823] =  'sd23800;
    data[7824] = -'sd44841;
    data[7825] = -'sd60364;
    data[7826] =  'sd25862;
    data[7827] = -'sd34531;
    data[7828] = -'sd8814;
    data[7829] = -'sd44070;
    data[7830] = -'sd56509;
    data[7831] =  'sd45137;
    data[7832] =  'sd61844;
    data[7833] = -'sd18462;
    data[7834] =  'sd71531;
    data[7835] =  'sd29973;
    data[7836] = -'sd13976;
    data[7837] = -'sd69880;
    data[7838] = -'sd21718;
    data[7839] =  'sd55251;
    data[7840] = -'sd51427;
    data[7841] =  'sd70547;
    data[7842] =  'sd25053;
    data[7843] = -'sd38576;
    data[7844] = -'sd29039;
    data[7845] =  'sd18646;
    data[7846] = -'sd70611;
    data[7847] = -'sd25373;
    data[7848] =  'sd36976;
    data[7849] =  'sd21039;
    data[7850] = -'sd58646;
    data[7851] =  'sd34452;
    data[7852] =  'sd8419;
    data[7853] =  'sd42095;
    data[7854] =  'sd46634;
    data[7855] =  'sd69329;
    data[7856] =  'sd18963;
    data[7857] = -'sd69026;
    data[7858] = -'sd17448;
    data[7859] =  'sd76601;
    data[7860] =  'sd55323;
    data[7861] = -'sd51067;
    data[7862] =  'sd72347;
    data[7863] =  'sd34053;
    data[7864] =  'sd6424;
    data[7865] =  'sd32120;
    data[7866] = -'sd3241;
    data[7867] = -'sd16205;
    data[7868] = -'sd81025;
    data[7869] = -'sd77443;
    data[7870] = -'sd59533;
    data[7871] =  'sd30017;
    data[7872] = -'sd13756;
    data[7873] = -'sd68780;
    data[7874] = -'sd16218;
    data[7875] = -'sd81090;
    data[7876] = -'sd77768;
    data[7877] = -'sd61158;
    data[7878] =  'sd21892;
    data[7879] = -'sd54381;
    data[7880] =  'sd55777;
    data[7881] = -'sd48797;
    data[7882] = -'sd80144;
    data[7883] = -'sd73038;
    data[7884] = -'sd37508;
    data[7885] = -'sd23699;
    data[7886] =  'sd45346;
    data[7887] =  'sd62889;
    data[7888] = -'sd13237;
    data[7889] = -'sd66185;
    data[7890] = -'sd3243;
    data[7891] = -'sd16215;
    data[7892] = -'sd81075;
    data[7893] = -'sd77693;
    data[7894] = -'sd60783;
    data[7895] =  'sd23767;
    data[7896] = -'sd45006;
    data[7897] = -'sd61189;
    data[7898] =  'sd21737;
    data[7899] = -'sd55156;
    data[7900] =  'sd51902;
    data[7901] = -'sd68172;
    data[7902] = -'sd13178;
    data[7903] = -'sd65890;
    data[7904] = -'sd1768;
    data[7905] = -'sd8840;
    data[7906] = -'sd44200;
    data[7907] = -'sd57159;
    data[7908] =  'sd41887;
    data[7909] =  'sd45594;
    data[7910] =  'sd64129;
    data[7911] = -'sd7037;
    data[7912] = -'sd35185;
    data[7913] = -'sd12084;
    data[7914] = -'sd60420;
    data[7915] =  'sd25582;
    data[7916] = -'sd35931;
    data[7917] = -'sd15814;
    data[7918] = -'sd79070;
    data[7919] = -'sd67668;
    data[7920] = -'sd10658;
    data[7921] = -'sd53290;
    data[7922] =  'sd61232;
    data[7923] = -'sd21522;
    data[7924] =  'sd56231;
    data[7925] = -'sd46527;
    data[7926] = -'sd68794;
    data[7927] = -'sd16288;
    data[7928] = -'sd81440;
    data[7929] = -'sd79518;
    data[7930] = -'sd69908;
    data[7931] = -'sd21858;
    data[7932] =  'sd54551;
    data[7933] = -'sd54927;
    data[7934] =  'sd53047;
    data[7935] = -'sd62447;
    data[7936] =  'sd15447;
    data[7937] =  'sd77235;
    data[7938] =  'sd58493;
    data[7939] = -'sd35217;
    data[7940] = -'sd12244;
    data[7941] = -'sd61220;
    data[7942] =  'sd21582;
    data[7943] = -'sd55931;
    data[7944] =  'sd48027;
    data[7945] =  'sd76294;
    data[7946] =  'sd53788;
    data[7947] = -'sd58742;
    data[7948] =  'sd33972;
    data[7949] =  'sd6019;
    data[7950] =  'sd30095;
    data[7951] = -'sd13366;
    data[7952] = -'sd66830;
    data[7953] = -'sd6468;
    data[7954] = -'sd32340;
    data[7955] =  'sd2141;
    data[7956] =  'sd10705;
    data[7957] =  'sd53525;
    data[7958] = -'sd60057;
    data[7959] =  'sd27397;
    data[7960] = -'sd26856;
    data[7961] =  'sd29561;
    data[7962] = -'sd16036;
    data[7963] = -'sd80180;
    data[7964] = -'sd73218;
    data[7965] = -'sd38408;
    data[7966] = -'sd28199;
    data[7967] =  'sd22846;
    data[7968] = -'sd49611;
    data[7969] =  'sd79627;
    data[7970] =  'sd70453;
    data[7971] =  'sd24583;
    data[7972] = -'sd40926;
    data[7973] = -'sd40789;
    data[7974] = -'sd40104;
    data[7975] = -'sd36679;
    data[7976] = -'sd19554;
    data[7977] =  'sd66071;
    data[7978] =  'sd2673;
    data[7979] =  'sd13365;
    data[7980] =  'sd66825;
    data[7981] =  'sd6443;
    data[7982] =  'sd32215;
    data[7983] = -'sd2766;
    data[7984] = -'sd13830;
    data[7985] = -'sd69150;
    data[7986] = -'sd18068;
    data[7987] =  'sd73501;
    data[7988] =  'sd39823;
    data[7989] =  'sd35274;
    data[7990] =  'sd12529;
    data[7991] =  'sd62645;
    data[7992] = -'sd14457;
    data[7993] = -'sd72285;
    data[7994] = -'sd33743;
    data[7995] = -'sd4874;
    data[7996] = -'sd24370;
    data[7997] =  'sd41991;
    data[7998] =  'sd46114;
    data[7999] =  'sd66729;
    data[8000] =  'sd5963;
    data[8001] =  'sd29815;
    data[8002] = -'sd14766;
    data[8003] = -'sd73830;
    data[8004] = -'sd41468;
    data[8005] = -'sd43499;
    data[8006] = -'sd53654;
    data[8007] =  'sd59412;
    data[8008] = -'sd30622;
    data[8009] =  'sd10731;
    data[8010] =  'sd53655;
    data[8011] = -'sd59407;
    data[8012] =  'sd30647;
    data[8013] = -'sd10606;
    data[8014] = -'sd53030;
    data[8015] =  'sd62532;
    data[8016] = -'sd15022;
    data[8017] = -'sd75110;
    data[8018] = -'sd47868;
    data[8019] = -'sd75499;
    data[8020] = -'sd49813;
    data[8021] =  'sd78617;
    data[8022] =  'sd65403;
    data[8023] = -'sd667;
    data[8024] = -'sd3335;
    data[8025] = -'sd16675;
    data[8026] =  'sd80466;
    data[8027] =  'sd74648;
    data[8028] =  'sd45558;
    data[8029] =  'sd63949;
    data[8030] = -'sd7937;
    data[8031] = -'sd39685;
    data[8032] = -'sd34584;
    data[8033] = -'sd9079;
    data[8034] = -'sd45395;
    data[8035] = -'sd63134;
    data[8036] =  'sd12012;
    data[8037] =  'sd60060;
    data[8038] = -'sd27382;
    data[8039] =  'sd26931;
    data[8040] = -'sd29186;
    data[8041] =  'sd17911;
    data[8042] = -'sd74286;
    data[8043] = -'sd43748;
    data[8044] = -'sd54899;
    data[8045] =  'sd53187;
    data[8046] = -'sd61747;
    data[8047] =  'sd18947;
    data[8048] = -'sd69106;
    data[8049] = -'sd17848;
    data[8050] =  'sd74601;
    data[8051] =  'sd45323;
    data[8052] =  'sd62774;
    data[8053] = -'sd13812;
    data[8054] = -'sd69060;
    data[8055] = -'sd17618;
    data[8056] =  'sd75751;
    data[8057] =  'sd51073;
    data[8058] = -'sd72317;
    data[8059] = -'sd33903;
    data[8060] = -'sd5674;
    data[8061] = -'sd28370;
    data[8062] =  'sd21991;
    data[8063] = -'sd53886;
    data[8064] =  'sd58252;
    data[8065] = -'sd36422;
    data[8066] = -'sd18269;
    data[8067] =  'sd72496;
    data[8068] =  'sd34798;
    data[8069] =  'sd10149;
    data[8070] =  'sd50745;
    data[8071] = -'sd73957;
    data[8072] = -'sd42103;
    data[8073] = -'sd46674;
    data[8074] = -'sd69529;
    data[8075] = -'sd19963;
    data[8076] =  'sd64026;
    data[8077] = -'sd7552;
    data[8078] = -'sd37760;
    data[8079] = -'sd24959;
    data[8080] =  'sd39046;
    data[8081] =  'sd31389;
    data[8082] = -'sd6896;
    data[8083] = -'sd34480;
    data[8084] = -'sd8559;
    data[8085] = -'sd42795;
    data[8086] = -'sd50134;
    data[8087] =  'sd77012;
    data[8088] =  'sd57378;
    data[8089] = -'sd40792;
    data[8090] = -'sd40119;
    data[8091] = -'sd36754;
    data[8092] = -'sd19929;
    data[8093] =  'sd64196;
    data[8094] = -'sd6702;
    data[8095] = -'sd33510;
    data[8096] = -'sd3709;
    data[8097] = -'sd18545;
    data[8098] =  'sd71116;
    data[8099] =  'sd27898;
    data[8100] = -'sd24351;
    data[8101] =  'sd42086;
    data[8102] =  'sd46589;
    data[8103] =  'sd69104;
    data[8104] =  'sd17838;
    data[8105] = -'sd74651;
    data[8106] = -'sd45573;
    data[8107] = -'sd64024;
    data[8108] =  'sd7562;
    data[8109] =  'sd37810;
    data[8110] =  'sd25209;
    data[8111] = -'sd37796;
    data[8112] = -'sd25139;
    data[8113] =  'sd38146;
    data[8114] =  'sd26889;
    data[8115] = -'sd29396;
    data[8116] =  'sd16861;
    data[8117] = -'sd79536;
    data[8118] = -'sd69998;
    data[8119] = -'sd22308;
    data[8120] =  'sd52301;
    data[8121] = -'sd66177;
    data[8122] = -'sd3203;
    data[8123] = -'sd16015;
    data[8124] = -'sd80075;
    data[8125] = -'sd72693;
    data[8126] = -'sd35783;
    data[8127] = -'sd15074;
    data[8128] = -'sd75370;
    data[8129] = -'sd49168;
    data[8130] =  'sd81842;
    data[8131] =  'sd81528;
    data[8132] =  'sd79958;
    data[8133] =  'sd72108;
    data[8134] =  'sd32858;
    data[8135] =  'sd449;
    data[8136] =  'sd2245;
    data[8137] =  'sd11225;
    data[8138] =  'sd56125;
    data[8139] = -'sd47057;
    data[8140] = -'sd71444;
    data[8141] = -'sd29538;
    data[8142] =  'sd16151;
    data[8143] =  'sd80755;
    data[8144] =  'sd76093;
    data[8145] =  'sd52783;
    data[8146] = -'sd63767;
    data[8147] =  'sd8847;
    data[8148] =  'sd44235;
    data[8149] =  'sd57334;
    data[8150] = -'sd41012;
    data[8151] = -'sd41219;
    data[8152] = -'sd42254;
    data[8153] = -'sd47429;
    data[8154] = -'sd73304;
    data[8155] = -'sd38838;
    data[8156] = -'sd30349;
    data[8157] =  'sd12096;
    data[8158] =  'sd60480;
    data[8159] = -'sd25282;
    data[8160] =  'sd37431;
    data[8161] =  'sd23314;
    data[8162] = -'sd47271;
    data[8163] = -'sd72514;
    data[8164] = -'sd34888;
    data[8165] = -'sd10599;
    data[8166] = -'sd52995;
    data[8167] =  'sd62707;
    data[8168] = -'sd14147;
    data[8169] = -'sd70735;
    data[8170] = -'sd25993;
    data[8171] =  'sd33876;
    data[8172] =  'sd5539;
    data[8173] =  'sd27695;
    data[8174] = -'sd25366;
    data[8175] =  'sd37011;
    data[8176] =  'sd21214;
    data[8177] = -'sd57771;
    data[8178] =  'sd38827;
    data[8179] =  'sd30294;
    data[8180] = -'sd12371;
    data[8181] = -'sd61855;
    data[8182] =  'sd18407;
    data[8183] = -'sd71806;
    data[8184] = -'sd31348;
    data[8185] =  'sd7101;
    data[8186] =  'sd35505;
    data[8187] =  'sd13684;
    data[8188] =  'sd68420;
    data[8189] =  'sd14418;
    data[8190] =  'sd72090;
    data[8191] =  'sd32768;
  end

endmodule

