module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd953;
  localparam R_DEPTH = 'd10;
  localparam B_LEN = 'd1505;
  localparam B_DEPTH = 'd11;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [13: 0] in_data;
  input      [10: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 14'h0f03; // 'd3843
      10'd1    : in_data <= 14'h056e; // 'd1390
      10'd2    : in_data <= 14'h0504; // 'd1284
      10'd3    : in_data <= 14'h0c49; // 'd3145
      10'd4    : in_data <= 14'h0b8c; // 'd2956
      10'd5    : in_data <= 14'h1738; // 'd5944
      10'd6    : in_data <= 14'h0dac; // 'd3500
      10'd7    : in_data <= 14'h0633; // 'd1587
      10'd8    : in_data <= 14'h11a1; // 'd4513
      10'd9    : in_data <= 14'h04ed; // 'd1261
      10'd10   : in_data <= 14'h0b76; // 'd2934
      10'd11   : in_data <= 14'h0de7; // 'd3559
      10'd12   : in_data <= 14'h007e; // 'd126
      10'd13   : in_data <= 14'h0d57; // 'd3415
      10'd14   : in_data <= 14'h1582; // 'd5506
      10'd15   : in_data <= 14'h0aab; // 'd2731
      10'd16   : in_data <= 14'h0f2b; // 'd3883
      10'd17   : in_data <= 14'h01e5; // 'd485
      10'd18   : in_data <= 14'h058d; // 'd1421
      10'd19   : in_data <= 14'h0698; // 'd1688
      10'd20   : in_data <= 14'h04b5; // 'd1205
      10'd21   : in_data <= 14'h0ecb; // 'd3787
      10'd22   : in_data <= 14'h15ce; // 'd5582
      10'd23   : in_data <= 14'h031e; // 'd798
      10'd24   : in_data <= 14'h0e81; // 'd3713
      10'd25   : in_data <= 14'h0677; // 'd1655
      10'd26   : in_data <= 14'h0ba2; // 'd2978
      10'd27   : in_data <= 14'h02bd; // 'd701
      10'd28   : in_data <= 14'h0606; // 'd1542
      10'd29   : in_data <= 14'h0302; // 'd770
      10'd30   : in_data <= 14'h0d62; // 'd3426
      10'd31   : in_data <= 14'h0301; // 'd769
      10'd32   : in_data <= 14'h01a3; // 'd419
      10'd33   : in_data <= 14'h063c; // 'd1596
      10'd34   : in_data <= 14'h0c9c; // 'd3228
      10'd35   : in_data <= 14'h161d; // 'd5661
      10'd36   : in_data <= 14'h0926; // 'd2342
      10'd37   : in_data <= 14'h1267; // 'd4711
      10'd38   : in_data <= 14'h00d2; // 'd210
      10'd39   : in_data <= 14'h096e; // 'd2414
      10'd40   : in_data <= 14'h0e79; // 'd3705
      10'd41   : in_data <= 14'h17bd; // 'd6077
      10'd42   : in_data <= 14'h169e; // 'd5790
      10'd43   : in_data <= 14'h0faf; // 'd4015
      10'd44   : in_data <= 14'h1625; // 'd5669
      10'd45   : in_data <= 14'h0b08; // 'd2824
      10'd46   : in_data <= 14'h0b18; // 'd2840
      10'd47   : in_data <= 14'h0631; // 'd1585
      10'd48   : in_data <= 14'h0dbf; // 'd3519
      10'd49   : in_data <= 14'h0538; // 'd1336
      10'd50   : in_data <= 14'h0d32; // 'd3378
      10'd51   : in_data <= 14'h1433; // 'd5171
      10'd52   : in_data <= 14'h0749; // 'd1865
      10'd53   : in_data <= 14'h111d; // 'd4381
      10'd54   : in_data <= 14'h02ff; // 'd767
      10'd55   : in_data <= 14'h0cfd; // 'd3325
      10'd56   : in_data <= 14'h120e; // 'd4622
      10'd57   : in_data <= 14'h0c85; // 'd3205
      10'd58   : in_data <= 14'h1122; // 'd4386
      10'd59   : in_data <= 14'h0414; // 'd1044
      10'd60   : in_data <= 14'h01c3; // 'd451
      10'd61   : in_data <= 14'h0b04; // 'd2820
      10'd62   : in_data <= 14'h04da; // 'd1242
      10'd63   : in_data <= 14'h0ae3; // 'd2787
      10'd64   : in_data <= 14'h1764; // 'd5988
      10'd65   : in_data <= 14'h0d59; // 'd3417
      10'd66   : in_data <= 14'h024b; // 'd587
      10'd67   : in_data <= 14'h0fea; // 'd4074
      10'd68   : in_data <= 14'h0b62; // 'd2914
      10'd69   : in_data <= 14'h16e5; // 'd5861
      10'd70   : in_data <= 14'h0efe; // 'd3838
      10'd71   : in_data <= 14'h00ad; // 'd173
      10'd72   : in_data <= 14'h0067; // 'd103
      10'd73   : in_data <= 14'h0c70; // 'd3184
      10'd74   : in_data <= 14'h0bc0; // 'd3008
      10'd75   : in_data <= 14'h1517; // 'd5399
      10'd76   : in_data <= 14'h10ef; // 'd4335
      10'd77   : in_data <= 14'h148b; // 'd5259
      10'd78   : in_data <= 14'h03f4; // 'd1012
      10'd79   : in_data <= 14'h092e; // 'd2350
      10'd80   : in_data <= 14'h0122; // 'd290
      10'd81   : in_data <= 14'h04de; // 'd1246
      10'd82   : in_data <= 14'h166f; // 'd5743
      10'd83   : in_data <= 14'h02b3; // 'd691
      10'd84   : in_data <= 14'h1131; // 'd4401
      10'd85   : in_data <= 14'h0264; // 'd612
      10'd86   : in_data <= 14'h08c3; // 'd2243
      10'd87   : in_data <= 14'h0f1e; // 'd3870
      10'd88   : in_data <= 14'h0d43; // 'd3395
      10'd89   : in_data <= 14'h14dc; // 'd5340
      10'd90   : in_data <= 14'h1514; // 'd5396
      10'd91   : in_data <= 14'h08ca; // 'd2250
      10'd92   : in_data <= 14'h13b1; // 'd5041
      10'd93   : in_data <= 14'h0d9c; // 'd3484
      10'd94   : in_data <= 14'h0946; // 'd2374
      10'd95   : in_data <= 14'h11fc; // 'd4604
      10'd96   : in_data <= 14'h18a6; // 'd6310
      10'd97   : in_data <= 14'h0bf9; // 'd3065
      10'd98   : in_data <= 14'h130e; // 'd4878
      10'd99   : in_data <= 14'h124a; // 'd4682
      10'd100  : in_data <= 14'h0cff; // 'd3327
      10'd101  : in_data <= 14'h12c0; // 'd4800
      10'd102  : in_data <= 14'h0675; // 'd1653
      10'd103  : in_data <= 14'h0f42; // 'd3906
      10'd104  : in_data <= 14'h0301; // 'd769
      10'd105  : in_data <= 14'h0940; // 'd2368
      10'd106  : in_data <= 14'h02e0; // 'd736
      10'd107  : in_data <= 14'h1093; // 'd4243
      10'd108  : in_data <= 14'h11f4; // 'd4596
      10'd109  : in_data <= 14'h0351; // 'd849
      10'd110  : in_data <= 14'h1891; // 'd6289
      10'd111  : in_data <= 14'h14bd; // 'd5309
      10'd112  : in_data <= 14'h0989; // 'd2441
      10'd113  : in_data <= 14'h0b1e; // 'd2846
      10'd114  : in_data <= 14'h1581; // 'd5505
      10'd115  : in_data <= 14'h0a6d; // 'd2669
      10'd116  : in_data <= 14'h1715; // 'd5909
      10'd117  : in_data <= 14'h138a; // 'd5002
      10'd118  : in_data <= 14'h0992; // 'd2450
      10'd119  : in_data <= 14'h1065; // 'd4197
      10'd120  : in_data <= 14'h0c98; // 'd3224
      10'd121  : in_data <= 14'h0d1e; // 'd3358
      10'd122  : in_data <= 14'h1748; // 'd5960
      10'd123  : in_data <= 14'h061d; // 'd1565
      10'd124  : in_data <= 14'h089b; // 'd2203
      10'd125  : in_data <= 14'h12e9; // 'd4841
      10'd126  : in_data <= 14'h00f7; // 'd247
      10'd127  : in_data <= 14'h035b; // 'd859
      10'd128  : in_data <= 14'h068e; // 'd1678
      10'd129  : in_data <= 14'h0007; // 'd7
      10'd130  : in_data <= 14'h0cf0; // 'd3312
      10'd131  : in_data <= 14'h03f0; // 'd1008
      10'd132  : in_data <= 14'h06fd; // 'd1789
      10'd133  : in_data <= 14'h0184; // 'd388
      10'd134  : in_data <= 14'h00b5; // 'd181
      10'd135  : in_data <= 14'h10d2; // 'd4306
      10'd136  : in_data <= 14'h0aa3; // 'd2723
      10'd137  : in_data <= 14'h1294; // 'd4756
      10'd138  : in_data <= 14'h11c8; // 'd4552
      10'd139  : in_data <= 14'h1891; // 'd6289
      10'd140  : in_data <= 14'h02cb; // 'd715
      10'd141  : in_data <= 14'h106a; // 'd4202
      10'd142  : in_data <= 14'h0f74; // 'd3956
      10'd143  : in_data <= 14'h1662; // 'd5730
      10'd144  : in_data <= 14'h0a0a; // 'd2570
      10'd145  : in_data <= 14'h0bd8; // 'd3032
      10'd146  : in_data <= 14'h16f2; // 'd5874
      10'd147  : in_data <= 14'h07b3; // 'd1971
      10'd148  : in_data <= 14'h0765; // 'd1893
      10'd149  : in_data <= 14'h050a; // 'd1290
      10'd150  : in_data <= 14'h0344; // 'd836
      10'd151  : in_data <= 14'h0fce; // 'd4046
      10'd152  : in_data <= 14'h0e86; // 'd3718
      10'd153  : in_data <= 14'h0278; // 'd632
      10'd154  : in_data <= 14'h07c1; // 'd1985
      10'd155  : in_data <= 14'h00d5; // 'd213
      10'd156  : in_data <= 14'h17d7; // 'd6103
      10'd157  : in_data <= 14'h12d0; // 'd4816
      10'd158  : in_data <= 14'h1089; // 'd4233
      10'd159  : in_data <= 14'h0a6d; // 'd2669
      10'd160  : in_data <= 14'h0f79; // 'd3961
      10'd161  : in_data <= 14'h0ca7; // 'd3239
      10'd162  : in_data <= 14'h01ae; // 'd430
      10'd163  : in_data <= 14'h12fa; // 'd4858
      10'd164  : in_data <= 14'h0311; // 'd785
      10'd165  : in_data <= 14'h0f13; // 'd3859
      10'd166  : in_data <= 14'h0336; // 'd822
      10'd167  : in_data <= 14'h0438; // 'd1080
      10'd168  : in_data <= 14'h0449; // 'd1097
      10'd169  : in_data <= 14'h05d8; // 'd1496
      10'd170  : in_data <= 14'h0a45; // 'd2629
      10'd171  : in_data <= 14'h0237; // 'd567
      10'd172  : in_data <= 14'h0008; // 'd8
      10'd173  : in_data <= 14'h189d; // 'd6301
      10'd174  : in_data <= 14'h0474; // 'd1140
      10'd175  : in_data <= 14'h1494; // 'd5268
      10'd176  : in_data <= 14'h0de1; // 'd3553
      10'd177  : in_data <= 14'h077c; // 'd1916
      10'd178  : in_data <= 14'h0a8d; // 'd2701
      10'd179  : in_data <= 14'h0b13; // 'd2835
      10'd180  : in_data <= 14'h05de; // 'd1502
      10'd181  : in_data <= 14'h1865; // 'd6245
      10'd182  : in_data <= 14'h05b9; // 'd1465
      10'd183  : in_data <= 14'h083a; // 'd2106
      10'd184  : in_data <= 14'h143c; // 'd5180
      10'd185  : in_data <= 14'h03f1; // 'd1009
      10'd186  : in_data <= 14'h09a4; // 'd2468
      10'd187  : in_data <= 14'h08d1; // 'd2257
      10'd188  : in_data <= 14'h00a2; // 'd162
      10'd189  : in_data <= 14'h1747; // 'd5959
      10'd190  : in_data <= 14'h09b6; // 'd2486
      10'd191  : in_data <= 14'h17c7; // 'd6087
      10'd192  : in_data <= 14'h03bd; // 'd957
      10'd193  : in_data <= 14'h163c; // 'd5692
      10'd194  : in_data <= 14'h015e; // 'd350
      10'd195  : in_data <= 14'h03fc; // 'd1020
      10'd196  : in_data <= 14'h17ed; // 'd6125
      10'd197  : in_data <= 14'h02da; // 'd730
      10'd198  : in_data <= 14'h1694; // 'd5780
      10'd199  : in_data <= 14'h09d0; // 'd2512
      10'd200  : in_data <= 14'h0436; // 'd1078
      10'd201  : in_data <= 14'h084e; // 'd2126
      10'd202  : in_data <= 14'h129e; // 'd4766
      10'd203  : in_data <= 14'h109e; // 'd4254
      10'd204  : in_data <= 14'h097b; // 'd2427
      10'd205  : in_data <= 14'h167e; // 'd5758
      10'd206  : in_data <= 14'h06a7; // 'd1703
      10'd207  : in_data <= 14'h1254; // 'd4692
      10'd208  : in_data <= 14'h12f3; // 'd4851
      10'd209  : in_data <= 14'h15b3; // 'd5555
      10'd210  : in_data <= 14'h17a0; // 'd6048
      10'd211  : in_data <= 14'h0b50; // 'd2896
      10'd212  : in_data <= 14'h046f; // 'd1135
      10'd213  : in_data <= 14'h06ae; // 'd1710
      10'd214  : in_data <= 14'h006b; // 'd107
      10'd215  : in_data <= 14'h0004; // 'd4
      10'd216  : in_data <= 14'h1836; // 'd6198
      10'd217  : in_data <= 14'h11f5; // 'd4597
      10'd218  : in_data <= 14'h0f5e; // 'd3934
      10'd219  : in_data <= 14'h0b46; // 'd2886
      10'd220  : in_data <= 14'h040b; // 'd1035
      10'd221  : in_data <= 14'h0ce8; // 'd3304
      10'd222  : in_data <= 14'h1893; // 'd6291
      10'd223  : in_data <= 14'h083f; // 'd2111
      10'd224  : in_data <= 14'h0586; // 'd1414
      10'd225  : in_data <= 14'h019d; // 'd413
      10'd226  : in_data <= 14'h0695; // 'd1685
      10'd227  : in_data <= 14'h13a6; // 'd5030
      10'd228  : in_data <= 14'h07f6; // 'd2038
      10'd229  : in_data <= 14'h098e; // 'd2446
      10'd230  : in_data <= 14'h0f43; // 'd3907
      10'd231  : in_data <= 14'h11f8; // 'd4600
      10'd232  : in_data <= 14'h05b4; // 'd1460
      10'd233  : in_data <= 14'h0897; // 'd2199
      10'd234  : in_data <= 14'h11e0; // 'd4576
      10'd235  : in_data <= 14'h02ab; // 'd683
      10'd236  : in_data <= 14'h1032; // 'd4146
      10'd237  : in_data <= 14'h06b3; // 'd1715
      10'd238  : in_data <= 14'h17f1; // 'd6129
      10'd239  : in_data <= 14'h0b15; // 'd2837
      10'd240  : in_data <= 14'h18b4; // 'd6324
      10'd241  : in_data <= 14'h16fe; // 'd5886
      10'd242  : in_data <= 14'h1124; // 'd4388
      10'd243  : in_data <= 14'h15cd; // 'd5581
      10'd244  : in_data <= 14'h143f; // 'd5183
      10'd245  : in_data <= 14'h0de7; // 'd3559
      10'd246  : in_data <= 14'h0920; // 'd2336
      10'd247  : in_data <= 14'h17e6; // 'd6118
      10'd248  : in_data <= 14'h17f5; // 'd6133
      10'd249  : in_data <= 14'h17ed; // 'd6125
      10'd250  : in_data <= 14'h16c6; // 'd5830
      10'd251  : in_data <= 14'h01ff; // 'd511
      10'd252  : in_data <= 14'h130b; // 'd4875
      10'd253  : in_data <= 14'h0fd1; // 'd4049
      10'd254  : in_data <= 14'h10df; // 'd4319
      10'd255  : in_data <= 14'h08c2; // 'd2242
      10'd256  : in_data <= 14'h145d; // 'd5213
      10'd257  : in_data <= 14'h07aa; // 'd1962
      10'd258  : in_data <= 14'h11fe; // 'd4606
      10'd259  : in_data <= 14'h06a6; // 'd1702
      10'd260  : in_data <= 14'h139b; // 'd5019
      10'd261  : in_data <= 14'h066e; // 'd1646
      10'd262  : in_data <= 14'h1029; // 'd4137
      10'd263  : in_data <= 14'h0e07; // 'd3591
      10'd264  : in_data <= 14'h1255; // 'd4693
      10'd265  : in_data <= 14'h07dc; // 'd2012
      10'd266  : in_data <= 14'h1223; // 'd4643
      10'd267  : in_data <= 14'h01c9; // 'd457
      10'd268  : in_data <= 14'h11b8; // 'd4536
      10'd269  : in_data <= 14'h0991; // 'd2449
      10'd270  : in_data <= 14'h02a6; // 'd678
      10'd271  : in_data <= 14'h0c56; // 'd3158
      10'd272  : in_data <= 14'h0c2d; // 'd3117
      10'd273  : in_data <= 14'h03e1; // 'd993
      10'd274  : in_data <= 14'h09a3; // 'd2467
      10'd275  : in_data <= 14'h0864; // 'd2148
      10'd276  : in_data <= 14'h0643; // 'd1603
      10'd277  : in_data <= 14'h11b1; // 'd4529
      10'd278  : in_data <= 14'h0f5f; // 'd3935
      10'd279  : in_data <= 14'h0949; // 'd2377
      10'd280  : in_data <= 14'h1684; // 'd5764
      10'd281  : in_data <= 14'h085f; // 'd2143
      10'd282  : in_data <= 14'h0941; // 'd2369
      10'd283  : in_data <= 14'h0e31; // 'd3633
      10'd284  : in_data <= 14'h145b; // 'd5211
      10'd285  : in_data <= 14'h015a; // 'd346
      10'd286  : in_data <= 14'h14f3; // 'd5363
      10'd287  : in_data <= 14'h0803; // 'd2051
      10'd288  : in_data <= 14'h127f; // 'd4735
      10'd289  : in_data <= 14'h0e07; // 'd3591
      10'd290  : in_data <= 14'h0860; // 'd2144
      10'd291  : in_data <= 14'h0eb0; // 'd3760
      10'd292  : in_data <= 14'h0f4c; // 'd3916
      10'd293  : in_data <= 14'h0f2f; // 'd3887
      10'd294  : in_data <= 14'h0548; // 'd1352
      10'd295  : in_data <= 14'h1152; // 'd4434
      10'd296  : in_data <= 14'h0e6f; // 'd3695
      10'd297  : in_data <= 14'h006f; // 'd111
      10'd298  : in_data <= 14'h025d; // 'd605
      10'd299  : in_data <= 14'h034a; // 'd842
      10'd300  : in_data <= 14'h1513; // 'd5395
      10'd301  : in_data <= 14'h0dd3; // 'd3539
      10'd302  : in_data <= 14'h0af0; // 'd2800
      10'd303  : in_data <= 14'h0763; // 'd1891
      10'd304  : in_data <= 14'h0894; // 'd2196
      10'd305  : in_data <= 14'h114e; // 'd4430
      10'd306  : in_data <= 14'h165b; // 'd5723
      10'd307  : in_data <= 14'h0723; // 'd1827
      10'd308  : in_data <= 14'h0f24; // 'd3876
      10'd309  : in_data <= 14'h1330; // 'd4912
      10'd310  : in_data <= 14'h0e6e; // 'd3694
      10'd311  : in_data <= 14'h0748; // 'd1864
      10'd312  : in_data <= 14'h155a; // 'd5466
      10'd313  : in_data <= 14'h18b8; // 'd6328
      10'd314  : in_data <= 14'h0985; // 'd2437
      10'd315  : in_data <= 14'h1435; // 'd5173
      10'd316  : in_data <= 14'h1285; // 'd4741
      10'd317  : in_data <= 14'h0578; // 'd1400
      10'd318  : in_data <= 14'h0532; // 'd1330
      10'd319  : in_data <= 14'h1898; // 'd6296
      10'd320  : in_data <= 14'h0c1a; // 'd3098
      10'd321  : in_data <= 14'h0366; // 'd870
      10'd322  : in_data <= 14'h0451; // 'd1105
      10'd323  : in_data <= 14'h16bb; // 'd5819
      10'd324  : in_data <= 14'h02f7; // 'd759
      10'd325  : in_data <= 14'h0703; // 'd1795
      10'd326  : in_data <= 14'h0db5; // 'd3509
      10'd327  : in_data <= 14'h13c6; // 'd5062
      10'd328  : in_data <= 14'h1144; // 'd4420
      10'd329  : in_data <= 14'h15d5; // 'd5589
      10'd330  : in_data <= 14'h077b; // 'd1915
      10'd331  : in_data <= 14'h16c0; // 'd5824
      10'd332  : in_data <= 14'h0c8b; // 'd3211
      10'd333  : in_data <= 14'h0545; // 'd1349
      10'd334  : in_data <= 14'h169b; // 'd5787
      10'd335  : in_data <= 14'h0264; // 'd612
      10'd336  : in_data <= 14'h08a6; // 'd2214
      10'd337  : in_data <= 14'h0d26; // 'd3366
      10'd338  : in_data <= 14'h0e07; // 'd3591
      10'd339  : in_data <= 14'h0e0b; // 'd3595
      10'd340  : in_data <= 14'h044b; // 'd1099
      10'd341  : in_data <= 14'h0204; // 'd516
      10'd342  : in_data <= 14'h12b2; // 'd4786
      10'd343  : in_data <= 14'h0b98; // 'd2968
      10'd344  : in_data <= 14'h0872; // 'd2162
      10'd345  : in_data <= 14'h0fac; // 'd4012
      10'd346  : in_data <= 14'h074f; // 'd1871
      10'd347  : in_data <= 14'h0eb5; // 'd3765
      10'd348  : in_data <= 14'h0ef5; // 'd3829
      10'd349  : in_data <= 14'h0467; // 'd1127
      10'd350  : in_data <= 14'h053f; // 'd1343
      10'd351  : in_data <= 14'h14cc; // 'd5324
      10'd352  : in_data <= 14'h08c5; // 'd2245
      10'd353  : in_data <= 14'h0ce6; // 'd3302
      10'd354  : in_data <= 14'h10ef; // 'd4335
      10'd355  : in_data <= 14'h0275; // 'd629
      10'd356  : in_data <= 14'h1427; // 'd5159
      10'd357  : in_data <= 14'h1242; // 'd4674
      10'd358  : in_data <= 14'h0098; // 'd152
      10'd359  : in_data <= 14'h031e; // 'd798
      10'd360  : in_data <= 14'h0131; // 'd305
      10'd361  : in_data <= 14'h03c4; // 'd964
      10'd362  : in_data <= 14'h04f7; // 'd1271
      10'd363  : in_data <= 14'h1800; // 'd6144
      10'd364  : in_data <= 14'h1182; // 'd4482
      10'd365  : in_data <= 14'h0d19; // 'd3353
      10'd366  : in_data <= 14'h0312; // 'd786
      10'd367  : in_data <= 14'h03a9; // 'd937
      10'd368  : in_data <= 14'h16c3; // 'd5827
      10'd369  : in_data <= 14'h0eb7; // 'd3767
      10'd370  : in_data <= 14'h0c48; // 'd3144
      10'd371  : in_data <= 14'h094a; // 'd2378
      10'd372  : in_data <= 14'h1829; // 'd6185
      10'd373  : in_data <= 14'h0d69; // 'd3433
      10'd374  : in_data <= 14'h02d4; // 'd724
      10'd375  : in_data <= 14'h02f1; // 'd753
      10'd376  : in_data <= 14'h1088; // 'd4232
      10'd377  : in_data <= 14'h0850; // 'd2128
      10'd378  : in_data <= 14'h1395; // 'd5013
      10'd379  : in_data <= 14'h0b3e; // 'd2878
      10'd380  : in_data <= 14'h02a4; // 'd676
      10'd381  : in_data <= 14'h00cb; // 'd203
      10'd382  : in_data <= 14'h09c9; // 'd2505
      10'd383  : in_data <= 14'h1832; // 'd6194
      10'd384  : in_data <= 14'h0caf; // 'd3247
      10'd385  : in_data <= 14'h0c82; // 'd3202
      10'd386  : in_data <= 14'h0d45; // 'd3397
      10'd387  : in_data <= 14'h14ad; // 'd5293
      10'd388  : in_data <= 14'h173c; // 'd5948
      10'd389  : in_data <= 14'h170e; // 'd5902
      10'd390  : in_data <= 14'h1039; // 'd4153
      10'd391  : in_data <= 14'h13d2; // 'd5074
      10'd392  : in_data <= 14'h0841; // 'd2113
      10'd393  : in_data <= 14'h0f32; // 'd3890
      10'd394  : in_data <= 14'h0dd5; // 'd3541
      10'd395  : in_data <= 14'h05a9; // 'd1449
      10'd396  : in_data <= 14'h0e0f; // 'd3599
      10'd397  : in_data <= 14'h018a; // 'd394
      10'd398  : in_data <= 14'h0788; // 'd1928
      10'd399  : in_data <= 14'h0a60; // 'd2656
      10'd400  : in_data <= 14'h10f3; // 'd4339
      10'd401  : in_data <= 14'h0145; // 'd325
      10'd402  : in_data <= 14'h15f5; // 'd5621
      10'd403  : in_data <= 14'h1465; // 'd5221
      10'd404  : in_data <= 14'h0879; // 'd2169
      10'd405  : in_data <= 14'h0725; // 'd1829
      10'd406  : in_data <= 14'h09f8; // 'd2552
      10'd407  : in_data <= 14'h00c4; // 'd196
      10'd408  : in_data <= 14'h0aa5; // 'd2725
      10'd409  : in_data <= 14'h1193; // 'd4499
      10'd410  : in_data <= 14'h0e9b; // 'd3739
      10'd411  : in_data <= 14'h0db8; // 'd3512
      10'd412  : in_data <= 14'h13b6; // 'd5046
      10'd413  : in_data <= 14'h088d; // 'd2189
      10'd414  : in_data <= 14'h0fcc; // 'd4044
      10'd415  : in_data <= 14'h0651; // 'd1617
      10'd416  : in_data <= 14'h15f0; // 'd5616
      10'd417  : in_data <= 14'h0b0e; // 'd2830
      10'd418  : in_data <= 14'h0173; // 'd371
      10'd419  : in_data <= 14'h127e; // 'd4734
      10'd420  : in_data <= 14'h17dd; // 'd6109
      10'd421  : in_data <= 14'h1052; // 'd4178
      10'd422  : in_data <= 14'h087f; // 'd2175
      10'd423  : in_data <= 14'h08a6; // 'd2214
      10'd424  : in_data <= 14'h0a23; // 'd2595
      10'd425  : in_data <= 14'h0dd7; // 'd3543
      10'd426  : in_data <= 14'h0dfa; // 'd3578
      10'd427  : in_data <= 14'h04b9; // 'd1209
      10'd428  : in_data <= 14'h1657; // 'd5719
      10'd429  : in_data <= 14'h0cd0; // 'd3280
      10'd430  : in_data <= 14'h03a0; // 'd928
      10'd431  : in_data <= 14'h0493; // 'd1171
      10'd432  : in_data <= 14'h0563; // 'd1379
      10'd433  : in_data <= 14'h0161; // 'd353
      10'd434  : in_data <= 14'h08f1; // 'd2289
      10'd435  : in_data <= 14'h061b; // 'd1563
      10'd436  : in_data <= 14'h0358; // 'd856
      10'd437  : in_data <= 14'h1532; // 'd5426
      10'd438  : in_data <= 14'h1520; // 'd5408
      10'd439  : in_data <= 14'h0d29; // 'd3369
      10'd440  : in_data <= 14'h15e0; // 'd5600
      10'd441  : in_data <= 14'h15d6; // 'd5590
      10'd442  : in_data <= 14'h0df9; // 'd3577
      10'd443  : in_data <= 14'h0034; // 'd52
      10'd444  : in_data <= 14'h1456; // 'd5206
      10'd445  : in_data <= 14'h0cc3; // 'd3267
      10'd446  : in_data <= 14'h01ad; // 'd429
      10'd447  : in_data <= 14'h1507; // 'd5383
      10'd448  : in_data <= 14'h0c79; // 'd3193
      10'd449  : in_data <= 14'h0c5e; // 'd3166
      10'd450  : in_data <= 14'h0769; // 'd1897
      10'd451  : in_data <= 14'h161e; // 'd5662
      10'd452  : in_data <= 14'h16de; // 'd5854
      10'd453  : in_data <= 14'h12a7; // 'd4775
      10'd454  : in_data <= 14'h0d19; // 'd3353
      10'd455  : in_data <= 14'h02d6; // 'd726
      10'd456  : in_data <= 14'h0364; // 'd868
      10'd457  : in_data <= 14'h11f1; // 'd4593
      10'd458  : in_data <= 14'h1225; // 'd4645
      10'd459  : in_data <= 14'h00d7; // 'd215
      10'd460  : in_data <= 14'h09af; // 'd2479
      10'd461  : in_data <= 14'h08b3; // 'd2227
      10'd462  : in_data <= 14'h0214; // 'd532
      10'd463  : in_data <= 14'h10b1; // 'd4273
      10'd464  : in_data <= 14'h10c4; // 'd4292
      10'd465  : in_data <= 14'h0cf9; // 'd3321
      10'd466  : in_data <= 14'h0c01; // 'd3073
      10'd467  : in_data <= 14'h13e5; // 'd5093
      10'd468  : in_data <= 14'h103f; // 'd4159
      10'd469  : in_data <= 14'h17a2; // 'd6050
      10'd470  : in_data <= 14'h00f2; // 'd242
      10'd471  : in_data <= 14'h0401; // 'd1025
      10'd472  : in_data <= 14'h1428; // 'd5160
      10'd473  : in_data <= 14'h0a0e; // 'd2574
      10'd474  : in_data <= 14'h0e61; // 'd3681
      10'd475  : in_data <= 14'h15f2; // 'd5618
      10'd476  : in_data <= 14'h162d; // 'd5677
      10'd477  : in_data <= 14'h013d; // 'd317
      10'd478  : in_data <= 14'h07d4; // 'd2004
      10'd479  : in_data <= 14'h0dfe; // 'd3582
      10'd480  : in_data <= 14'h1382; // 'd4994
      10'd481  : in_data <= 14'h06c2; // 'd1730
      10'd482  : in_data <= 14'h12a7; // 'd4775
      10'd483  : in_data <= 14'h07df; // 'd2015
      10'd484  : in_data <= 14'h035c; // 'd860
      10'd485  : in_data <= 14'h1486; // 'd5254
      10'd486  : in_data <= 14'h15cb; // 'd5579
      10'd487  : in_data <= 14'h06d5; // 'd1749
      10'd488  : in_data <= 14'h0e3f; // 'd3647
      10'd489  : in_data <= 14'h05bb; // 'd1467
      10'd490  : in_data <= 14'h16e1; // 'd5857
      10'd491  : in_data <= 14'h0f0b; // 'd3851
      10'd492  : in_data <= 14'h0d18; // 'd3352
      10'd493  : in_data <= 14'h109c; // 'd4252
      10'd494  : in_data <= 14'h08cc; // 'd2252
      10'd495  : in_data <= 14'h0ac8; // 'd2760
      10'd496  : in_data <= 14'h0ee2; // 'd3810
      10'd497  : in_data <= 14'h0dee; // 'd3566
      10'd498  : in_data <= 14'h1812; // 'd6162
      10'd499  : in_data <= 14'h0d27; // 'd3367
      10'd500  : in_data <= 14'h01fb; // 'd507
      10'd501  : in_data <= 14'h0068; // 'd104
      10'd502  : in_data <= 14'h0315; // 'd789
      10'd503  : in_data <= 14'h0933; // 'd2355
      10'd504  : in_data <= 14'h06fa; // 'd1786
      10'd505  : in_data <= 14'h0f44; // 'd3908
      10'd506  : in_data <= 14'h0117; // 'd279
      10'd507  : in_data <= 14'h057d; // 'd1405
      10'd508  : in_data <= 14'h171d; // 'd5917
      10'd509  : in_data <= 14'h072b; // 'd1835
      10'd510  : in_data <= 14'h0802; // 'd2050
      10'd511  : in_data <= 14'h165a; // 'd5722
      10'd512  : in_data <= 14'h02c5; // 'd709
      10'd513  : in_data <= 14'h0ee8; // 'd3816
      10'd514  : in_data <= 14'h0c0b; // 'd3083
      10'd515  : in_data <= 14'h0e25; // 'd3621
      10'd516  : in_data <= 14'h01ca; // 'd458
      10'd517  : in_data <= 14'h0239; // 'd569
      10'd518  : in_data <= 14'h1607; // 'd5639
      10'd519  : in_data <= 14'h0011; // 'd17
      10'd520  : in_data <= 14'h0aee; // 'd2798
      10'd521  : in_data <= 14'h0613; // 'd1555
      10'd522  : in_data <= 14'h1893; // 'd6291
      10'd523  : in_data <= 14'h0d8a; // 'd3466
      10'd524  : in_data <= 14'h1451; // 'd5201
      10'd525  : in_data <= 14'h0282; // 'd642
      10'd526  : in_data <= 14'h0f2b; // 'd3883
      10'd527  : in_data <= 14'h0501; // 'd1281
      10'd528  : in_data <= 14'h04a4; // 'd1188
      10'd529  : in_data <= 14'h1655; // 'd5717
      10'd530  : in_data <= 14'h010c; // 'd268
      10'd531  : in_data <= 14'h06ae; // 'd1710
      10'd532  : in_data <= 14'h12b0; // 'd4784
      10'd533  : in_data <= 14'h1282; // 'd4738
      10'd534  : in_data <= 14'h007f; // 'd127
      10'd535  : in_data <= 14'h15cc; // 'd5580
      10'd536  : in_data <= 14'h069a; // 'd1690
      10'd537  : in_data <= 14'h01b1; // 'd433
      10'd538  : in_data <= 14'h0857; // 'd2135
      10'd539  : in_data <= 14'h153a; // 'd5434
      10'd540  : in_data <= 14'h0b73; // 'd2931
      10'd541  : in_data <= 14'h07fe; // 'd2046
      10'd542  : in_data <= 14'h07f5; // 'd2037
      10'd543  : in_data <= 14'h0cdc; // 'd3292
      10'd544  : in_data <= 14'h08a5; // 'd2213
      10'd545  : in_data <= 14'h1226; // 'd4646
      10'd546  : in_data <= 14'h1197; // 'd4503
      10'd547  : in_data <= 14'h10bf; // 'd4287
      10'd548  : in_data <= 14'h0c14; // 'd3092
      10'd549  : in_data <= 14'h11b9; // 'd4537
      10'd550  : in_data <= 14'h098f; // 'd2447
      10'd551  : in_data <= 14'h1641; // 'd5697
      10'd552  : in_data <= 14'h0eed; // 'd3821
      10'd553  : in_data <= 14'h0294; // 'd660
      10'd554  : in_data <= 14'h089b; // 'd2203
      10'd555  : in_data <= 14'h16a9; // 'd5801
      10'd556  : in_data <= 14'h06d8; // 'd1752
      10'd557  : in_data <= 14'h03e8; // 'd1000
      10'd558  : in_data <= 14'h0ce7; // 'd3303
      10'd559  : in_data <= 14'h1399; // 'd5017
      10'd560  : in_data <= 14'h0dd4; // 'd3540
      10'd561  : in_data <= 14'h0071; // 'd113
      10'd562  : in_data <= 14'h11a0; // 'd4512
      10'd563  : in_data <= 14'h0da5; // 'd3493
      10'd564  : in_data <= 14'h0d61; // 'd3425
      10'd565  : in_data <= 14'h0caa; // 'd3242
      10'd566  : in_data <= 14'h00c0; // 'd192
      10'd567  : in_data <= 14'h107d; // 'd4221
      10'd568  : in_data <= 14'h17bb; // 'd6075
      10'd569  : in_data <= 14'h03f7; // 'd1015
      10'd570  : in_data <= 14'h1670; // 'd5744
      10'd571  : in_data <= 14'h1767; // 'd5991
      10'd572  : in_data <= 14'h1258; // 'd4696
      10'd573  : in_data <= 14'h165a; // 'd5722
      10'd574  : in_data <= 14'h0808; // 'd2056
      10'd575  : in_data <= 14'h179e; // 'd6046
      10'd576  : in_data <= 14'h009e; // 'd158
      10'd577  : in_data <= 14'h146b; // 'd5227
      10'd578  : in_data <= 14'h0e22; // 'd3618
      10'd579  : in_data <= 14'h0570; // 'd1392
      10'd580  : in_data <= 14'h15e6; // 'd5606
      10'd581  : in_data <= 14'h08de; // 'd2270
      10'd582  : in_data <= 14'h0188; // 'd392
      10'd583  : in_data <= 14'h10f1; // 'd4337
      10'd584  : in_data <= 14'h0aa1; // 'd2721
      10'd585  : in_data <= 14'h04fc; // 'd1276
      10'd586  : in_data <= 14'h021a; // 'd538
      10'd587  : in_data <= 14'h1787; // 'd6023
      10'd588  : in_data <= 14'h11cc; // 'd4556
      10'd589  : in_data <= 14'h1187; // 'd4487
      10'd590  : in_data <= 14'h1814; // 'd6164
      10'd591  : in_data <= 14'h0b32; // 'd2866
      10'd592  : in_data <= 14'h10f3; // 'd4339
      10'd593  : in_data <= 14'h12e9; // 'd4841
      10'd594  : in_data <= 14'h08c6; // 'd2246
      10'd595  : in_data <= 14'h11cc; // 'd4556
      10'd596  : in_data <= 14'h065c; // 'd1628
      10'd597  : in_data <= 14'h17dc; // 'd6108
      10'd598  : in_data <= 14'h044f; // 'd1103
      10'd599  : in_data <= 14'h166b; // 'd5739
      10'd600  : in_data <= 14'h1365; // 'd4965
      10'd601  : in_data <= 14'h05fc; // 'd1532
      10'd602  : in_data <= 14'h10bc; // 'd4284
      10'd603  : in_data <= 14'h01b1; // 'd433
      10'd604  : in_data <= 14'h0ea2; // 'd3746
      10'd605  : in_data <= 14'h10a9; // 'd4265
      10'd606  : in_data <= 14'h1471; // 'd5233
      10'd607  : in_data <= 14'h09a4; // 'd2468
      10'd608  : in_data <= 14'h0526; // 'd1318
      10'd609  : in_data <= 14'h175d; // 'd5981
      10'd610  : in_data <= 14'h0812; // 'd2066
      10'd611  : in_data <= 14'h0f62; // 'd3938
      10'd612  : in_data <= 14'h1019; // 'd4121
      10'd613  : in_data <= 14'h00ae; // 'd174
      10'd614  : in_data <= 14'h11a9; // 'd4521
      10'd615  : in_data <= 14'h074d; // 'd1869
      10'd616  : in_data <= 14'h1174; // 'd4468
      10'd617  : in_data <= 14'h16c9; // 'd5833
      10'd618  : in_data <= 14'h13de; // 'd5086
      10'd619  : in_data <= 14'h162d; // 'd5677
      10'd620  : in_data <= 14'h1607; // 'd5639
      10'd621  : in_data <= 14'h0365; // 'd869
      10'd622  : in_data <= 14'h0be1; // 'd3041
      10'd623  : in_data <= 14'h0dc8; // 'd3528
      10'd624  : in_data <= 14'h0e22; // 'd3618
      10'd625  : in_data <= 14'h0191; // 'd401
      10'd626  : in_data <= 14'h103c; // 'd4156
      10'd627  : in_data <= 14'h0e6f; // 'd3695
      10'd628  : in_data <= 14'h163b; // 'd5691
      10'd629  : in_data <= 14'h136a; // 'd4970
      10'd630  : in_data <= 14'h0e27; // 'd3623
      10'd631  : in_data <= 14'h0604; // 'd1540
      10'd632  : in_data <= 14'h018e; // 'd398
      10'd633  : in_data <= 14'h143e; // 'd5182
      10'd634  : in_data <= 14'h0a7d; // 'd2685
      10'd635  : in_data <= 14'h0787; // 'd1927
      10'd636  : in_data <= 14'h136a; // 'd4970
      10'd637  : in_data <= 14'h0f33; // 'd3891
      10'd638  : in_data <= 14'h085e; // 'd2142
      10'd639  : in_data <= 14'h03b2; // 'd946
      10'd640  : in_data <= 14'h11b7; // 'd4535
      10'd641  : in_data <= 14'h16d6; // 'd5846
      10'd642  : in_data <= 14'h0747; // 'd1863
      10'd643  : in_data <= 14'h129d; // 'd4765
      10'd644  : in_data <= 14'h15c1; // 'd5569
      10'd645  : in_data <= 14'h1634; // 'd5684
      10'd646  : in_data <= 14'h05a8; // 'd1448
      10'd647  : in_data <= 14'h010a; // 'd266
      10'd648  : in_data <= 14'h0d21; // 'd3361
      10'd649  : in_data <= 14'h17dc; // 'd6108
      10'd650  : in_data <= 14'h02d5; // 'd725
      10'd651  : in_data <= 14'h049e; // 'd1182
      10'd652  : in_data <= 14'h1676; // 'd5750
      10'd653  : in_data <= 14'h160f; // 'd5647
      10'd654  : in_data <= 14'h10da; // 'd4314
      10'd655  : in_data <= 14'h127e; // 'd4734
      10'd656  : in_data <= 14'h1386; // 'd4998
      10'd657  : in_data <= 14'h03a0; // 'd928
      10'd658  : in_data <= 14'h0d3b; // 'd3387
      10'd659  : in_data <= 14'h0afd; // 'd2813
      10'd660  : in_data <= 14'h0d5f; // 'd3423
      10'd661  : in_data <= 14'h107a; // 'd4218
      10'd662  : in_data <= 14'h04f8; // 'd1272
      10'd663  : in_data <= 14'h0316; // 'd790
      10'd664  : in_data <= 14'h13df; // 'd5087
      10'd665  : in_data <= 14'h0009; // 'd9
      10'd666  : in_data <= 14'h017e; // 'd382
      10'd667  : in_data <= 14'h02b6; // 'd694
      10'd668  : in_data <= 14'h01cc; // 'd460
      10'd669  : in_data <= 14'h13bf; // 'd5055
      10'd670  : in_data <= 14'h0a01; // 'd2561
      10'd671  : in_data <= 14'h132a; // 'd4906
      10'd672  : in_data <= 14'h07c5; // 'd1989
      10'd673  : in_data <= 14'h0a06; // 'd2566
      10'd674  : in_data <= 14'h1782; // 'd6018
      10'd675  : in_data <= 14'h0a24; // 'd2596
      10'd676  : in_data <= 14'h09bf; // 'd2495
      10'd677  : in_data <= 14'h00be; // 'd190
      10'd678  : in_data <= 14'h0357; // 'd855
      10'd679  : in_data <= 14'h173d; // 'd5949
      10'd680  : in_data <= 14'h0d53; // 'd3411
      10'd681  : in_data <= 14'h0ecc; // 'd3788
      10'd682  : in_data <= 14'h081e; // 'd2078
      10'd683  : in_data <= 14'h118c; // 'd4492
      10'd684  : in_data <= 14'h146b; // 'd5227
      10'd685  : in_data <= 14'h127f; // 'd4735
      10'd686  : in_data <= 14'h1789; // 'd6025
      10'd687  : in_data <= 14'h0d78; // 'd3448
      10'd688  : in_data <= 14'h0b4e; // 'd2894
      10'd689  : in_data <= 14'h05bc; // 'd1468
      10'd690  : in_data <= 14'h09de; // 'd2526
      10'd691  : in_data <= 14'h0068; // 'd104
      10'd692  : in_data <= 14'h0d8b; // 'd3467
      10'd693  : in_data <= 14'h1138; // 'd4408
      10'd694  : in_data <= 14'h11c5; // 'd4549
      10'd695  : in_data <= 14'h06ac; // 'd1708
      10'd696  : in_data <= 14'h0b5c; // 'd2908
      10'd697  : in_data <= 14'h0ab6; // 'd2742
      10'd698  : in_data <= 14'h173d; // 'd5949
      10'd699  : in_data <= 14'h04fc; // 'd1276
      10'd700  : in_data <= 14'h0917; // 'd2327
      10'd701  : in_data <= 14'h1477; // 'd5239
      10'd702  : in_data <= 14'h13fc; // 'd5116
      10'd703  : in_data <= 14'h0633; // 'd1587
      10'd704  : in_data <= 14'h087b; // 'd2171
      10'd705  : in_data <= 14'h05ea; // 'd1514
      10'd706  : in_data <= 14'h11c8; // 'd4552
      10'd707  : in_data <= 14'h0547; // 'd1351
      10'd708  : in_data <= 14'h1787; // 'd6023
      10'd709  : in_data <= 14'h07dc; // 'd2012
      10'd710  : in_data <= 14'h1198; // 'd4504
      10'd711  : in_data <= 14'h05c4; // 'd1476
      10'd712  : in_data <= 14'h1374; // 'd4980
      10'd713  : in_data <= 14'h111e; // 'd4382
      10'd714  : in_data <= 14'h04f2; // 'd1266
      10'd715  : in_data <= 14'h0d32; // 'd3378
      10'd716  : in_data <= 14'h088d; // 'd2189
      10'd717  : in_data <= 14'h048c; // 'd1164
      10'd718  : in_data <= 14'h1005; // 'd4101
      10'd719  : in_data <= 14'h04a4; // 'd1188
      10'd720  : in_data <= 14'h0f8b; // 'd3979
      10'd721  : in_data <= 14'h171c; // 'd5916
      10'd722  : in_data <= 14'h0580; // 'd1408
      10'd723  : in_data <= 14'h0c7c; // 'd3196
      10'd724  : in_data <= 14'h02fc; // 'd764
      10'd725  : in_data <= 14'h0108; // 'd264
      10'd726  : in_data <= 14'h038f; // 'd911
      10'd727  : in_data <= 14'h0c4b; // 'd3147
      10'd728  : in_data <= 14'h0872; // 'd2162
      10'd729  : in_data <= 14'h14ce; // 'd5326
      10'd730  : in_data <= 14'h0f09; // 'd3849
      10'd731  : in_data <= 14'h16bd; // 'd5821
      10'd732  : in_data <= 14'h01eb; // 'd491
      10'd733  : in_data <= 14'h170e; // 'd5902
      10'd734  : in_data <= 14'h0533; // 'd1331
      10'd735  : in_data <= 14'h1647; // 'd5703
      10'd736  : in_data <= 14'h0b4a; // 'd2890
      10'd737  : in_data <= 14'h1497; // 'd5271
      10'd738  : in_data <= 14'h051a; // 'd1306
      10'd739  : in_data <= 14'h03d0; // 'd976
      10'd740  : in_data <= 14'h1346; // 'd4934
      10'd741  : in_data <= 14'h10a7; // 'd4263
      10'd742  : in_data <= 14'h1650; // 'd5712
      10'd743  : in_data <= 14'h041e; // 'd1054
      10'd744  : in_data <= 14'h0513; // 'd1299
      10'd745  : in_data <= 14'h0484; // 'd1156
      10'd746  : in_data <= 14'h0ba2; // 'd2978
      10'd747  : in_data <= 14'h16c4; // 'd5828
      10'd748  : in_data <= 14'h08ca; // 'd2250
      10'd749  : in_data <= 14'h000d; // 'd13
      10'd750  : in_data <= 14'h0728; // 'd1832
      10'd751  : in_data <= 14'h1253; // 'd4691
      10'd752  : in_data <= 14'h099c; // 'd2460
      10'd753  : in_data <= 14'h1696; // 'd5782
      10'd754  : in_data <= 14'h058c; // 'd1420
      10'd755  : in_data <= 14'h016d; // 'd365
      10'd756  : in_data <= 14'h048b; // 'd1163
      10'd757  : in_data <= 14'h0368; // 'd872
      10'd758  : in_data <= 14'h0230; // 'd560
      10'd759  : in_data <= 14'h0bd5; // 'd3029
      10'd760  : in_data <= 14'h163f; // 'd5695
      10'd761  : in_data <= 14'h05a3; // 'd1443
      10'd762  : in_data <= 14'h01cd; // 'd461
      10'd763  : in_data <= 14'h164f; // 'd5711
      10'd764  : in_data <= 14'h038f; // 'd911
      10'd765  : in_data <= 14'h0eab; // 'd3755
      10'd766  : in_data <= 14'h16cd; // 'd5837
      10'd767  : in_data <= 14'h123b; // 'd4667
      10'd768  : in_data <= 14'h02c6; // 'd710
      10'd769  : in_data <= 14'h09ad; // 'd2477
      10'd770  : in_data <= 14'h0378; // 'd888
      10'd771  : in_data <= 14'h15bb; // 'd5563
      10'd772  : in_data <= 14'h0587; // 'd1415
      10'd773  : in_data <= 14'h13cd; // 'd5069
      10'd774  : in_data <= 14'h034e; // 'd846
      10'd775  : in_data <= 14'h0b76; // 'd2934
      10'd776  : in_data <= 14'h16fd; // 'd5885
      10'd777  : in_data <= 14'h0c22; // 'd3106
      10'd778  : in_data <= 14'h0c09; // 'd3081
      10'd779  : in_data <= 14'h0cf6; // 'd3318
      10'd780  : in_data <= 14'h1326; // 'd4902
      10'd781  : in_data <= 14'h1735; // 'd5941
      10'd782  : in_data <= 14'h01b5; // 'd437
      10'd783  : in_data <= 14'h0a77; // 'd2679
      10'd784  : in_data <= 14'h12f4; // 'd4852
      10'd785  : in_data <= 14'h05f9; // 'd1529
      10'd786  : in_data <= 14'h11b1; // 'd4529
      10'd787  : in_data <= 14'h167f; // 'd5759
      10'd788  : in_data <= 14'h1768; // 'd5992
      10'd789  : in_data <= 14'h0b46; // 'd2886
      10'd790  : in_data <= 14'h0a28; // 'd2600
      10'd791  : in_data <= 14'h0d42; // 'd3394
      10'd792  : in_data <= 14'h045c; // 'd1116
      10'd793  : in_data <= 14'h17d3; // 'd6099
      10'd794  : in_data <= 14'h06fa; // 'd1786
      10'd795  : in_data <= 14'h1529; // 'd5417
      10'd796  : in_data <= 14'h0169; // 'd361
      10'd797  : in_data <= 14'h179f; // 'd6047
      10'd798  : in_data <= 14'h00fd; // 'd253
      10'd799  : in_data <= 14'h07aa; // 'd1962
      10'd800  : in_data <= 14'h0f90; // 'd3984
      10'd801  : in_data <= 14'h0681; // 'd1665
      10'd802  : in_data <= 14'h0331; // 'd817
      10'd803  : in_data <= 14'h15f6; // 'd5622
      10'd804  : in_data <= 14'h0aa2; // 'd2722
      10'd805  : in_data <= 14'h171e; // 'd5918
      10'd806  : in_data <= 14'h0de1; // 'd3553
      10'd807  : in_data <= 14'h1037; // 'd4151
      10'd808  : in_data <= 14'h066d; // 'd1645
      10'd809  : in_data <= 14'h0e2a; // 'd3626
      10'd810  : in_data <= 14'h1850; // 'd6224
      10'd811  : in_data <= 14'h137f; // 'd4991
      10'd812  : in_data <= 14'h0c20; // 'd3104
      10'd813  : in_data <= 14'h0902; // 'd2306
      10'd814  : in_data <= 14'h17c8; // 'd6088
      10'd815  : in_data <= 14'h0565; // 'd1381
      10'd816  : in_data <= 14'h11d6; // 'd4566
      10'd817  : in_data <= 14'h0edc; // 'd3804
      10'd818  : in_data <= 14'h04b8; // 'd1208
      10'd819  : in_data <= 14'h12ed; // 'd4845
      10'd820  : in_data <= 14'h1796; // 'd6038
      10'd821  : in_data <= 14'h03e4; // 'd996
      10'd822  : in_data <= 14'h0b18; // 'd2840
      10'd823  : in_data <= 14'h0ca8; // 'd3240
      10'd824  : in_data <= 14'h0a65; // 'd2661
      10'd825  : in_data <= 14'h0196; // 'd406
      10'd826  : in_data <= 14'h07eb; // 'd2027
      10'd827  : in_data <= 14'h0233; // 'd563
      10'd828  : in_data <= 14'h0670; // 'd1648
      10'd829  : in_data <= 14'h171b; // 'd5915
      10'd830  : in_data <= 14'h143a; // 'd5178
      10'd831  : in_data <= 14'h0363; // 'd867
      10'd832  : in_data <= 14'h1772; // 'd6002
      10'd833  : in_data <= 14'h0c85; // 'd3205
      10'd834  : in_data <= 14'h12ac; // 'd4780
      10'd835  : in_data <= 14'h10f9; // 'd4345
      10'd836  : in_data <= 14'h0bdf; // 'd3039
      10'd837  : in_data <= 14'h03f1; // 'd1009
      10'd838  : in_data <= 14'h0821; // 'd2081
      10'd839  : in_data <= 14'h0899; // 'd2201
      10'd840  : in_data <= 14'h11ba; // 'd4538
      10'd841  : in_data <= 14'h11af; // 'd4527
      10'd842  : in_data <= 14'h0d9c; // 'd3484
      10'd843  : in_data <= 14'h0086; // 'd134
      10'd844  : in_data <= 14'h12fd; // 'd4861
      10'd845  : in_data <= 14'h1123; // 'd4387
      10'd846  : in_data <= 14'h0335; // 'd821
      10'd847  : in_data <= 14'h07cd; // 'd1997
      10'd848  : in_data <= 14'h0ffe; // 'd4094
      10'd849  : in_data <= 14'h06bf; // 'd1727
      10'd850  : in_data <= 14'h13f6; // 'd5110
      10'd851  : in_data <= 14'h0db1; // 'd3505
      10'd852  : in_data <= 14'h0665; // 'd1637
      10'd853  : in_data <= 14'h09b8; // 'd2488
      10'd854  : in_data <= 14'h0d7c; // 'd3452
      10'd855  : in_data <= 14'h1435; // 'd5173
      10'd856  : in_data <= 14'h0daa; // 'd3498
      10'd857  : in_data <= 14'h106d; // 'd4205
      10'd858  : in_data <= 14'h1754; // 'd5972
      10'd859  : in_data <= 14'h0f20; // 'd3872
      10'd860  : in_data <= 14'h1400; // 'd5120
      10'd861  : in_data <= 14'h0e01; // 'd3585
      10'd862  : in_data <= 14'h15e1; // 'd5601
      10'd863  : in_data <= 14'h0a99; // 'd2713
      10'd864  : in_data <= 14'h0e39; // 'd3641
      10'd865  : in_data <= 14'h1888; // 'd6280
      10'd866  : in_data <= 14'h0b50; // 'd2896
      10'd867  : in_data <= 14'h0799; // 'd1945
      10'd868  : in_data <= 14'h113c; // 'd4412
      10'd869  : in_data <= 14'h1429; // 'd5161
      10'd870  : in_data <= 14'h0ac3; // 'd2755
      10'd871  : in_data <= 14'h0729; // 'd1833
      10'd872  : in_data <= 14'h13a5; // 'd5029
      10'd873  : in_data <= 14'h10dd; // 'd4317
      10'd874  : in_data <= 14'h0d59; // 'd3417
      10'd875  : in_data <= 14'h039a; // 'd922
      10'd876  : in_data <= 14'h175b; // 'd5979
      10'd877  : in_data <= 14'h067c; // 'd1660
      10'd878  : in_data <= 14'h07bb; // 'd1979
      10'd879  : in_data <= 14'h022a; // 'd554
      10'd880  : in_data <= 14'h01ad; // 'd429
      10'd881  : in_data <= 14'h1219; // 'd4633
      10'd882  : in_data <= 14'h0cc7; // 'd3271
      10'd883  : in_data <= 14'h0fb2; // 'd4018
      10'd884  : in_data <= 14'h14b8; // 'd5304
      10'd885  : in_data <= 14'h125a; // 'd4698
      10'd886  : in_data <= 14'h0845; // 'd2117
      10'd887  : in_data <= 14'h1399; // 'd5017
      10'd888  : in_data <= 14'h0638; // 'd1592
      10'd889  : in_data <= 14'h1754; // 'd5972
      10'd890  : in_data <= 14'h00a3; // 'd163
      10'd891  : in_data <= 14'h0e52; // 'd3666
      10'd892  : in_data <= 14'h0e00; // 'd3584
      10'd893  : in_data <= 14'h1169; // 'd4457
      10'd894  : in_data <= 14'h06c4; // 'd1732
      10'd895  : in_data <= 14'h171a; // 'd5914
      10'd896  : in_data <= 14'h14a7; // 'd5287
      10'd897  : in_data <= 14'h1348; // 'd4936
      10'd898  : in_data <= 14'h17eb; // 'd6123
      10'd899  : in_data <= 14'h0241; // 'd577
      10'd900  : in_data <= 14'h0655; // 'd1621
      10'd901  : in_data <= 14'h1653; // 'd5715
      10'd902  : in_data <= 14'h12d1; // 'd4817
      10'd903  : in_data <= 14'h02d8; // 'd728
      10'd904  : in_data <= 14'h1054; // 'd4180
      10'd905  : in_data <= 14'h0b35; // 'd2869
      10'd906  : in_data <= 14'h187d; // 'd6269
      10'd907  : in_data <= 14'h0a4e; // 'd2638
      10'd908  : in_data <= 14'h02dc; // 'd732
      10'd909  : in_data <= 14'h0ee2; // 'd3810
      10'd910  : in_data <= 14'h0bef; // 'd3055
      10'd911  : in_data <= 14'h172a; // 'd5930
      10'd912  : in_data <= 14'h007d; // 'd125
      10'd913  : in_data <= 14'h01ab; // 'd427
      10'd914  : in_data <= 14'h0caf; // 'd3247
      10'd915  : in_data <= 14'h0ba8; // 'd2984
      10'd916  : in_data <= 14'h0792; // 'd1938
      10'd917  : in_data <= 14'h11b8; // 'd4536
      10'd918  : in_data <= 14'h167e; // 'd5758
      10'd919  : in_data <= 14'h0c5f; // 'd3167
      10'd920  : in_data <= 14'h029f; // 'd671
      10'd921  : in_data <= 14'h0a8f; // 'd2703
      10'd922  : in_data <= 14'h052e; // 'd1326
      10'd923  : in_data <= 14'h18af; // 'd6319
      10'd924  : in_data <= 14'h04f0; // 'd1264
      10'd925  : in_data <= 14'h0fc4; // 'd4036
      10'd926  : in_data <= 14'h070b; // 'd1803
      10'd927  : in_data <= 14'h00a4; // 'd164
      10'd928  : in_data <= 14'h06e1; // 'd1761
      10'd929  : in_data <= 14'h10ed; // 'd4333
      10'd930  : in_data <= 14'h04af; // 'd1199
      10'd931  : in_data <= 14'h1568; // 'd5480
      10'd932  : in_data <= 14'h0ae9; // 'd2793
      10'd933  : in_data <= 14'h17d9; // 'd6105
      10'd934  : in_data <= 14'h10e9; // 'd4329
      10'd935  : in_data <= 14'h0d9c; // 'd3484
      10'd936  : in_data <= 14'h0d2f; // 'd3375
      10'd937  : in_data <= 14'h04d0; // 'd1232
      10'd938  : in_data <= 14'h10ee; // 'd4334
      10'd939  : in_data <= 14'h0213; // 'd531
      10'd940  : in_data <= 14'h15b5; // 'd5557
      10'd941  : in_data <= 14'h0474; // 'd1140
      10'd942  : in_data <= 14'h101d; // 'd4125
      10'd943  : in_data <= 14'h0a00; // 'd2560
      10'd944  : in_data <= 14'h14d5; // 'd5333
      10'd945  : in_data <= 14'h13a1; // 'd5025
      10'd946  : in_data <= 14'h1411; // 'd5137
      10'd947  : in_data <= 14'h1262; // 'd4706
      10'd948  : in_data <= 14'h0370; // 'd880
      10'd949  : in_data <= 14'h00ee; // 'd238
      10'd950  : in_data <= 14'h15e7; // 'd5607
      10'd951  : in_data <= 14'h18b2; // 'd6322
      10'd952  : in_data <= 14'h0c76; // 'd3190
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      11'd0    : out_data_ref <= 8'h85;
      11'd1    : out_data_ref <= 8'h97;
      11'd2    : out_data_ref <= 8'hc3;
      11'd3    : out_data_ref <= 8'h69;
      11'd4    : out_data_ref <= 8'h14;
      11'd5    : out_data_ref <= 8'h58;
      11'd6    : out_data_ref <= 8'h51;
      11'd7    : out_data_ref <= 8'ha7;
      11'd8    : out_data_ref <= 8'hdc;
      11'd9    : out_data_ref <= 8'h1d;
      11'd10   : out_data_ref <= 8'h07;
      11'd11   : out_data_ref <= 8'h82;
      11'd12   : out_data_ref <= 8'h1f;
      11'd13   : out_data_ref <= 8'h87;
      11'd14   : out_data_ref <= 8'h6f;
      11'd15   : out_data_ref <= 8'h68;
      11'd16   : out_data_ref <= 8'h2e;
      11'd17   : out_data_ref <= 8'h00;
      11'd18   : out_data_ref <= 8'hb5;
      11'd19   : out_data_ref <= 8'h65;
      11'd20   : out_data_ref <= 8'h82;
      11'd21   : out_data_ref <= 8'h8c;
      11'd22   : out_data_ref <= 8'h20;
      11'd23   : out_data_ref <= 8'h52;
      11'd24   : out_data_ref <= 8'h02;
      11'd25   : out_data_ref <= 8'h3d;
      11'd26   : out_data_ref <= 8'h8d;
      11'd27   : out_data_ref <= 8'he4;
      11'd28   : out_data_ref <= 8'h94;
      11'd29   : out_data_ref <= 8'h8c;
      11'd30   : out_data_ref <= 8'h29;
      11'd31   : out_data_ref <= 8'h7b;
      11'd32   : out_data_ref <= 8'h47;
      11'd33   : out_data_ref <= 8'h7a;
      11'd34   : out_data_ref <= 8'h27;
      11'd35   : out_data_ref <= 8'hf5;
      11'd36   : out_data_ref <= 8'h37;
      11'd37   : out_data_ref <= 8'hff;
      11'd38   : out_data_ref <= 8'h54;
      11'd39   : out_data_ref <= 8'ha5;
      11'd40   : out_data_ref <= 8'h64;
      11'd41   : out_data_ref <= 8'h3a;
      11'd42   : out_data_ref <= 8'ha7;
      11'd43   : out_data_ref <= 8'haf;
      11'd44   : out_data_ref <= 8'h5d;
      11'd45   : out_data_ref <= 8'h69;
      11'd46   : out_data_ref <= 8'h2f;
      11'd47   : out_data_ref <= 8'h73;
      11'd48   : out_data_ref <= 8'h47;
      11'd49   : out_data_ref <= 8'h5c;
      11'd50   : out_data_ref <= 8'hd7;
      11'd51   : out_data_ref <= 8'h88;
      11'd52   : out_data_ref <= 8'hd4;
      11'd53   : out_data_ref <= 8'h0c;
      11'd54   : out_data_ref <= 8'haa;
      11'd55   : out_data_ref <= 8'hd3;
      11'd56   : out_data_ref <= 8'h71;
      11'd57   : out_data_ref <= 8'h45;
      11'd58   : out_data_ref <= 8'hae;
      11'd59   : out_data_ref <= 8'h1c;
      11'd60   : out_data_ref <= 8'hdf;
      11'd61   : out_data_ref <= 8'hf1;
      11'd62   : out_data_ref <= 8'h4f;
      11'd63   : out_data_ref <= 8'hc3;
      11'd64   : out_data_ref <= 8'h93;
      11'd65   : out_data_ref <= 8'hcf;
      11'd66   : out_data_ref <= 8'h31;
      11'd67   : out_data_ref <= 8'h51;
      11'd68   : out_data_ref <= 8'h65;
      11'd69   : out_data_ref <= 8'h4f;
      11'd70   : out_data_ref <= 8'h79;
      11'd71   : out_data_ref <= 8'hcd;
      11'd72   : out_data_ref <= 8'h77;
      11'd73   : out_data_ref <= 8'h2b;
      11'd74   : out_data_ref <= 8'ha1;
      11'd75   : out_data_ref <= 8'h98;
      11'd76   : out_data_ref <= 8'hfc;
      11'd77   : out_data_ref <= 8'h10;
      11'd78   : out_data_ref <= 8'hb6;
      11'd79   : out_data_ref <= 8'h76;
      11'd80   : out_data_ref <= 8'hb4;
      11'd81   : out_data_ref <= 8'h99;
      11'd82   : out_data_ref <= 8'h94;
      11'd83   : out_data_ref <= 8'hf7;
      11'd84   : out_data_ref <= 8'hed;
      11'd85   : out_data_ref <= 8'h4c;
      11'd86   : out_data_ref <= 8'h15;
      11'd87   : out_data_ref <= 8'h99;
      11'd88   : out_data_ref <= 8'h47;
      11'd89   : out_data_ref <= 8'he4;
      11'd90   : out_data_ref <= 8'h1a;
      11'd91   : out_data_ref <= 8'hda;
      11'd92   : out_data_ref <= 8'hf5;
      11'd93   : out_data_ref <= 8'h47;
      11'd94   : out_data_ref <= 8'h2a;
      11'd95   : out_data_ref <= 8'ha4;
      11'd96   : out_data_ref <= 8'h35;
      11'd97   : out_data_ref <= 8'hbf;
      11'd98   : out_data_ref <= 8'h94;
      11'd99   : out_data_ref <= 8'h3a;
      11'd100  : out_data_ref <= 8'h3f;
      11'd101  : out_data_ref <= 8'ha0;
      11'd102  : out_data_ref <= 8'hc3;
      11'd103  : out_data_ref <= 8'h12;
      11'd104  : out_data_ref <= 8'hc1;
      11'd105  : out_data_ref <= 8'h33;
      11'd106  : out_data_ref <= 8'h25;
      11'd107  : out_data_ref <= 8'had;
      11'd108  : out_data_ref <= 8'heb;
      11'd109  : out_data_ref <= 8'h3d;
      11'd110  : out_data_ref <= 8'h7c;
      11'd111  : out_data_ref <= 8'hef;
      11'd112  : out_data_ref <= 8'hdb;
      11'd113  : out_data_ref <= 8'h7d;
      11'd114  : out_data_ref <= 8'h3c;
      11'd115  : out_data_ref <= 8'h68;
      11'd116  : out_data_ref <= 8'h5b;
      11'd117  : out_data_ref <= 8'h37;
      11'd118  : out_data_ref <= 8'h15;
      11'd119  : out_data_ref <= 8'h40;
      11'd120  : out_data_ref <= 8'hea;
      11'd121  : out_data_ref <= 8'h0e;
      11'd122  : out_data_ref <= 8'hd3;
      11'd123  : out_data_ref <= 8'h8f;
      11'd124  : out_data_ref <= 8'hba;
      11'd125  : out_data_ref <= 8'h93;
      11'd126  : out_data_ref <= 8'hb4;
      11'd127  : out_data_ref <= 8'h24;
      11'd128  : out_data_ref <= 8'hff;
      11'd129  : out_data_ref <= 8'hb3;
      11'd130  : out_data_ref <= 8'h80;
      11'd131  : out_data_ref <= 8'h9c;
      11'd132  : out_data_ref <= 8'h99;
      11'd133  : out_data_ref <= 8'h94;
      11'd134  : out_data_ref <= 8'hf3;
      11'd135  : out_data_ref <= 8'hc3;
      11'd136  : out_data_ref <= 8'haf;
      11'd137  : out_data_ref <= 8'h5b;
      11'd138  : out_data_ref <= 8'h7f;
      11'd139  : out_data_ref <= 8'hc2;
      11'd140  : out_data_ref <= 8'h31;
      11'd141  : out_data_ref <= 8'hb5;
      11'd142  : out_data_ref <= 8'ha2;
      11'd143  : out_data_ref <= 8'ha5;
      11'd144  : out_data_ref <= 8'hf2;
      11'd145  : out_data_ref <= 8'h7e;
      11'd146  : out_data_ref <= 8'h17;
      11'd147  : out_data_ref <= 8'hdb;
      11'd148  : out_data_ref <= 8'h2b;
      11'd149  : out_data_ref <= 8'he2;
      11'd150  : out_data_ref <= 8'h66;
      11'd151  : out_data_ref <= 8'h9c;
      11'd152  : out_data_ref <= 8'hce;
      11'd153  : out_data_ref <= 8'h39;
      11'd154  : out_data_ref <= 8'h54;
      11'd155  : out_data_ref <= 8'ha5;
      11'd156  : out_data_ref <= 8'h87;
      11'd157  : out_data_ref <= 8'h37;
      11'd158  : out_data_ref <= 8'h44;
      11'd159  : out_data_ref <= 8'h63;
      11'd160  : out_data_ref <= 8'h4a;
      11'd161  : out_data_ref <= 8'h8d;
      11'd162  : out_data_ref <= 8'h04;
      11'd163  : out_data_ref <= 8'h32;
      11'd164  : out_data_ref <= 8'hd6;
      11'd165  : out_data_ref <= 8'h82;
      11'd166  : out_data_ref <= 8'hbe;
      11'd167  : out_data_ref <= 8'h8a;
      11'd168  : out_data_ref <= 8'h31;
      11'd169  : out_data_ref <= 8'hcf;
      11'd170  : out_data_ref <= 8'h06;
      11'd171  : out_data_ref <= 8'heb;
      11'd172  : out_data_ref <= 8'h13;
      11'd173  : out_data_ref <= 8'hda;
      11'd174  : out_data_ref <= 8'h80;
      11'd175  : out_data_ref <= 8'he3;
      11'd176  : out_data_ref <= 8'h45;
      11'd177  : out_data_ref <= 8'h7f;
      11'd178  : out_data_ref <= 8'h52;
      11'd179  : out_data_ref <= 8'h6e;
      11'd180  : out_data_ref <= 8'h61;
      11'd181  : out_data_ref <= 8'h74;
      11'd182  : out_data_ref <= 8'hcf;
      11'd183  : out_data_ref <= 8'hda;
      11'd184  : out_data_ref <= 8'h93;
      11'd185  : out_data_ref <= 8'hbc;
      11'd186  : out_data_ref <= 8'h1b;
      11'd187  : out_data_ref <= 8'h7c;
      11'd188  : out_data_ref <= 8'hd3;
      11'd189  : out_data_ref <= 8'hc0;
      11'd190  : out_data_ref <= 8'h67;
      11'd191  : out_data_ref <= 8'h2d;
      11'd192  : out_data_ref <= 8'h61;
      11'd193  : out_data_ref <= 8'hec;
      11'd194  : out_data_ref <= 8'h42;
      11'd195  : out_data_ref <= 8'hba;
      11'd196  : out_data_ref <= 8'h63;
      11'd197  : out_data_ref <= 8'hbf;
      11'd198  : out_data_ref <= 8'h44;
      11'd199  : out_data_ref <= 8'h37;
      11'd200  : out_data_ref <= 8'hd8;
      11'd201  : out_data_ref <= 8'hc8;
      11'd202  : out_data_ref <= 8'h70;
      11'd203  : out_data_ref <= 8'hcd;
      11'd204  : out_data_ref <= 8'h6d;
      11'd205  : out_data_ref <= 8'h55;
      11'd206  : out_data_ref <= 8'hf3;
      11'd207  : out_data_ref <= 8'h25;
      11'd208  : out_data_ref <= 8'h18;
      11'd209  : out_data_ref <= 8'hb9;
      11'd210  : out_data_ref <= 8'hd0;
      11'd211  : out_data_ref <= 8'h62;
      11'd212  : out_data_ref <= 8'hb1;
      11'd213  : out_data_ref <= 8'h85;
      11'd214  : out_data_ref <= 8'h87;
      11'd215  : out_data_ref <= 8'h63;
      11'd216  : out_data_ref <= 8'ha9;
      11'd217  : out_data_ref <= 8'h05;
      11'd218  : out_data_ref <= 8'hc8;
      11'd219  : out_data_ref <= 8'h62;
      11'd220  : out_data_ref <= 8'h63;
      11'd221  : out_data_ref <= 8'hcc;
      11'd222  : out_data_ref <= 8'h8c;
      11'd223  : out_data_ref <= 8'h69;
      11'd224  : out_data_ref <= 8'h91;
      11'd225  : out_data_ref <= 8'hfe;
      11'd226  : out_data_ref <= 8'h9f;
      11'd227  : out_data_ref <= 8'hdc;
      11'd228  : out_data_ref <= 8'h58;
      11'd229  : out_data_ref <= 8'hc5;
      11'd230  : out_data_ref <= 8'h0b;
      11'd231  : out_data_ref <= 8'h47;
      11'd232  : out_data_ref <= 8'h15;
      11'd233  : out_data_ref <= 8'hdb;
      11'd234  : out_data_ref <= 8'hcd;
      11'd235  : out_data_ref <= 8'h2c;
      11'd236  : out_data_ref <= 8'h57;
      11'd237  : out_data_ref <= 8'h0d;
      11'd238  : out_data_ref <= 8'h44;
      11'd239  : out_data_ref <= 8'had;
      11'd240  : out_data_ref <= 8'h26;
      11'd241  : out_data_ref <= 8'hc8;
      11'd242  : out_data_ref <= 8'h7f;
      11'd243  : out_data_ref <= 8'h3b;
      11'd244  : out_data_ref <= 8'hd0;
      11'd245  : out_data_ref <= 8'h8a;
      11'd246  : out_data_ref <= 8'hea;
      11'd247  : out_data_ref <= 8'h2c;
      11'd248  : out_data_ref <= 8'h30;
      11'd249  : out_data_ref <= 8'he9;
      11'd250  : out_data_ref <= 8'hff;
      11'd251  : out_data_ref <= 8'h8b;
      11'd252  : out_data_ref <= 8'h82;
      11'd253  : out_data_ref <= 8'hf6;
      11'd254  : out_data_ref <= 8'had;
      11'd255  : out_data_ref <= 8'h0f;
      11'd256  : out_data_ref <= 8'h83;
      11'd257  : out_data_ref <= 8'hf9;
      11'd258  : out_data_ref <= 8'h08;
      11'd259  : out_data_ref <= 8'hcd;
      11'd260  : out_data_ref <= 8'h1d;
      11'd261  : out_data_ref <= 8'h63;
      11'd262  : out_data_ref <= 8'h9a;
      11'd263  : out_data_ref <= 8'h9f;
      11'd264  : out_data_ref <= 8'h59;
      11'd265  : out_data_ref <= 8'hce;
      11'd266  : out_data_ref <= 8'h62;
      11'd267  : out_data_ref <= 8'h4d;
      11'd268  : out_data_ref <= 8'h6f;
      11'd269  : out_data_ref <= 8'h19;
      11'd270  : out_data_ref <= 8'h80;
      11'd271  : out_data_ref <= 8'ha9;
      11'd272  : out_data_ref <= 8'h14;
      11'd273  : out_data_ref <= 8'h28;
      11'd274  : out_data_ref <= 8'h5f;
      11'd275  : out_data_ref <= 8'hef;
      11'd276  : out_data_ref <= 8'hda;
      11'd277  : out_data_ref <= 8'h5e;
      11'd278  : out_data_ref <= 8'h1e;
      11'd279  : out_data_ref <= 8'h1f;
      11'd280  : out_data_ref <= 8'h5d;
      11'd281  : out_data_ref <= 8'h80;
      11'd282  : out_data_ref <= 8'h58;
      11'd283  : out_data_ref <= 8'ha9;
      11'd284  : out_data_ref <= 8'h51;
      11'd285  : out_data_ref <= 8'h91;
      11'd286  : out_data_ref <= 8'h48;
      11'd287  : out_data_ref <= 8'h97;
      11'd288  : out_data_ref <= 8'hf0;
      11'd289  : out_data_ref <= 8'ha1;
      11'd290  : out_data_ref <= 8'h30;
      11'd291  : out_data_ref <= 8'hf3;
      11'd292  : out_data_ref <= 8'hd5;
      11'd293  : out_data_ref <= 8'h44;
      11'd294  : out_data_ref <= 8'h06;
      11'd295  : out_data_ref <= 8'h2c;
      11'd296  : out_data_ref <= 8'hb8;
      11'd297  : out_data_ref <= 8'hcc;
      11'd298  : out_data_ref <= 8'he3;
      11'd299  : out_data_ref <= 8'h80;
      11'd300  : out_data_ref <= 8'h18;
      11'd301  : out_data_ref <= 8'h9c;
      11'd302  : out_data_ref <= 8'he5;
      11'd303  : out_data_ref <= 8'h10;
      11'd304  : out_data_ref <= 8'h36;
      11'd305  : out_data_ref <= 8'hcc;
      11'd306  : out_data_ref <= 8'h90;
      11'd307  : out_data_ref <= 8'hea;
      11'd308  : out_data_ref <= 8'h74;
      11'd309  : out_data_ref <= 8'h79;
      11'd310  : out_data_ref <= 8'h66;
      11'd311  : out_data_ref <= 8'h77;
      11'd312  : out_data_ref <= 8'h62;
      11'd313  : out_data_ref <= 8'h8c;
      11'd314  : out_data_ref <= 8'hb8;
      11'd315  : out_data_ref <= 8'hb6;
      11'd316  : out_data_ref <= 8'hcd;
      11'd317  : out_data_ref <= 8'h92;
      11'd318  : out_data_ref <= 8'h5a;
      11'd319  : out_data_ref <= 8'h63;
      11'd320  : out_data_ref <= 8'h64;
      11'd321  : out_data_ref <= 8'h40;
      11'd322  : out_data_ref <= 8'hae;
      11'd323  : out_data_ref <= 8'h37;
      11'd324  : out_data_ref <= 8'h4c;
      11'd325  : out_data_ref <= 8'hbe;
      11'd326  : out_data_ref <= 8'h9f;
      11'd327  : out_data_ref <= 8'hfc;
      11'd328  : out_data_ref <= 8'hd7;
      11'd329  : out_data_ref <= 8'h01;
      11'd330  : out_data_ref <= 8'hbb;
      11'd331  : out_data_ref <= 8'hb6;
      11'd332  : out_data_ref <= 8'h2e;
      11'd333  : out_data_ref <= 8'h9d;
      11'd334  : out_data_ref <= 8'h57;
      11'd335  : out_data_ref <= 8'h52;
      11'd336  : out_data_ref <= 8'h30;
      11'd337  : out_data_ref <= 8'hd1;
      11'd338  : out_data_ref <= 8'h94;
      11'd339  : out_data_ref <= 8'h00;
      11'd340  : out_data_ref <= 8'h67;
      11'd341  : out_data_ref <= 8'hf5;
      11'd342  : out_data_ref <= 8'hda;
      11'd343  : out_data_ref <= 8'h55;
      11'd344  : out_data_ref <= 8'h26;
      11'd345  : out_data_ref <= 8'h57;
      11'd346  : out_data_ref <= 8'h02;
      11'd347  : out_data_ref <= 8'h6e;
      11'd348  : out_data_ref <= 8'h06;
      11'd349  : out_data_ref <= 8'h23;
      11'd350  : out_data_ref <= 8'hd3;
      11'd351  : out_data_ref <= 8'h4f;
      11'd352  : out_data_ref <= 8'h8f;
      11'd353  : out_data_ref <= 8'h9f;
      11'd354  : out_data_ref <= 8'he2;
      11'd355  : out_data_ref <= 8'hf1;
      11'd356  : out_data_ref <= 8'h75;
      11'd357  : out_data_ref <= 8'h75;
      11'd358  : out_data_ref <= 8'hea;
      11'd359  : out_data_ref <= 8'h3c;
      11'd360  : out_data_ref <= 8'h8d;
      11'd361  : out_data_ref <= 8'h4e;
      11'd362  : out_data_ref <= 8'hf7;
      11'd363  : out_data_ref <= 8'hac;
      11'd364  : out_data_ref <= 8'hf1;
      11'd365  : out_data_ref <= 8'h97;
      11'd366  : out_data_ref <= 8'h71;
      11'd367  : out_data_ref <= 8'hb3;
      11'd368  : out_data_ref <= 8'h04;
      11'd369  : out_data_ref <= 8'haf;
      11'd370  : out_data_ref <= 8'hce;
      11'd371  : out_data_ref <= 8'h34;
      11'd372  : out_data_ref <= 8'hc8;
      11'd373  : out_data_ref <= 8'h5c;
      11'd374  : out_data_ref <= 8'h2b;
      11'd375  : out_data_ref <= 8'he4;
      11'd376  : out_data_ref <= 8'hb8;
      11'd377  : out_data_ref <= 8'h06;
      11'd378  : out_data_ref <= 8'hc7;
      11'd379  : out_data_ref <= 8'ha0;
      11'd380  : out_data_ref <= 8'h71;
      11'd381  : out_data_ref <= 8'ha8;
      11'd382  : out_data_ref <= 8'ha7;
      11'd383  : out_data_ref <= 8'h88;
      11'd384  : out_data_ref <= 8'hbd;
      11'd385  : out_data_ref <= 8'hf5;
      11'd386  : out_data_ref <= 8'hc0;
      11'd387  : out_data_ref <= 8'h57;
      11'd388  : out_data_ref <= 8'h1e;
      11'd389  : out_data_ref <= 8'h53;
      11'd390  : out_data_ref <= 8'h77;
      11'd391  : out_data_ref <= 8'h28;
      11'd392  : out_data_ref <= 8'h1f;
      11'd393  : out_data_ref <= 8'h88;
      11'd394  : out_data_ref <= 8'h34;
      11'd395  : out_data_ref <= 8'h4c;
      11'd396  : out_data_ref <= 8'h55;
      11'd397  : out_data_ref <= 8'h30;
      11'd398  : out_data_ref <= 8'h28;
      11'd399  : out_data_ref <= 8'h18;
      11'd400  : out_data_ref <= 8'h96;
      11'd401  : out_data_ref <= 8'h85;
      11'd402  : out_data_ref <= 8'h78;
      11'd403  : out_data_ref <= 8'h68;
      11'd404  : out_data_ref <= 8'h3c;
      11'd405  : out_data_ref <= 8'h0e;
      11'd406  : out_data_ref <= 8'h54;
      11'd407  : out_data_ref <= 8'h02;
      11'd408  : out_data_ref <= 8'hea;
      11'd409  : out_data_ref <= 8'h7b;
      11'd410  : out_data_ref <= 8'ha3;
      11'd411  : out_data_ref <= 8'hf8;
      11'd412  : out_data_ref <= 8'h51;
      11'd413  : out_data_ref <= 8'hf1;
      11'd414  : out_data_ref <= 8'hc3;
      11'd415  : out_data_ref <= 8'h90;
      11'd416  : out_data_ref <= 8'hd2;
      11'd417  : out_data_ref <= 8'hfd;
      11'd418  : out_data_ref <= 8'h65;
      11'd419  : out_data_ref <= 8'h31;
      11'd420  : out_data_ref <= 8'h9b;
      11'd421  : out_data_ref <= 8'h77;
      11'd422  : out_data_ref <= 8'h89;
      11'd423  : out_data_ref <= 8'h51;
      11'd424  : out_data_ref <= 8'h44;
      11'd425  : out_data_ref <= 8'hf4;
      11'd426  : out_data_ref <= 8'hc9;
      11'd427  : out_data_ref <= 8'h11;
      11'd428  : out_data_ref <= 8'h07;
      11'd429  : out_data_ref <= 8'h8c;
      11'd430  : out_data_ref <= 8'he5;
      11'd431  : out_data_ref <= 8'h59;
      11'd432  : out_data_ref <= 8'hca;
      11'd433  : out_data_ref <= 8'h2f;
      11'd434  : out_data_ref <= 8'hee;
      11'd435  : out_data_ref <= 8'h4f;
      11'd436  : out_data_ref <= 8'h36;
      11'd437  : out_data_ref <= 8'h2d;
      11'd438  : out_data_ref <= 8'hff;
      11'd439  : out_data_ref <= 8'h27;
      11'd440  : out_data_ref <= 8'h3a;
      11'd441  : out_data_ref <= 8'h1f;
      11'd442  : out_data_ref <= 8'h65;
      11'd443  : out_data_ref <= 8'h16;
      11'd444  : out_data_ref <= 8'heb;
      11'd445  : out_data_ref <= 8'h47;
      11'd446  : out_data_ref <= 8'h1e;
      11'd447  : out_data_ref <= 8'h02;
      11'd448  : out_data_ref <= 8'h8b;
      11'd449  : out_data_ref <= 8'h79;
      11'd450  : out_data_ref <= 8'hbb;
      11'd451  : out_data_ref <= 8'h08;
      11'd452  : out_data_ref <= 8'haf;
      11'd453  : out_data_ref <= 8'h3e;
      11'd454  : out_data_ref <= 8'h73;
      11'd455  : out_data_ref <= 8'h51;
      11'd456  : out_data_ref <= 8'hbb;
      11'd457  : out_data_ref <= 8'h8d;
      11'd458  : out_data_ref <= 8'h46;
      11'd459  : out_data_ref <= 8'he1;
      11'd460  : out_data_ref <= 8'hd4;
      11'd461  : out_data_ref <= 8'h94;
      11'd462  : out_data_ref <= 8'hab;
      11'd463  : out_data_ref <= 8'h93;
      11'd464  : out_data_ref <= 8'h53;
      11'd465  : out_data_ref <= 8'h7e;
      11'd466  : out_data_ref <= 8'h04;
      11'd467  : out_data_ref <= 8'hfb;
      11'd468  : out_data_ref <= 8'h2d;
      11'd469  : out_data_ref <= 8'h9f;
      11'd470  : out_data_ref <= 8'hb9;
      11'd471  : out_data_ref <= 8'h35;
      11'd472  : out_data_ref <= 8'h0a;
      11'd473  : out_data_ref <= 8'h35;
      11'd474  : out_data_ref <= 8'h7f;
      11'd475  : out_data_ref <= 8'hcd;
      11'd476  : out_data_ref <= 8'h98;
      11'd477  : out_data_ref <= 8'hc4;
      11'd478  : out_data_ref <= 8'h46;
      11'd479  : out_data_ref <= 8'hb8;
      11'd480  : out_data_ref <= 8'h50;
      11'd481  : out_data_ref <= 8'h84;
      11'd482  : out_data_ref <= 8'h00;
      11'd483  : out_data_ref <= 8'h19;
      11'd484  : out_data_ref <= 8'h86;
      11'd485  : out_data_ref <= 8'h87;
      11'd486  : out_data_ref <= 8'h5e;
      11'd487  : out_data_ref <= 8'h5d;
      11'd488  : out_data_ref <= 8'h9c;
      11'd489  : out_data_ref <= 8'h0a;
      11'd490  : out_data_ref <= 8'h6e;
      11'd491  : out_data_ref <= 8'hd0;
      11'd492  : out_data_ref <= 8'h5c;
      11'd493  : out_data_ref <= 8'h96;
      11'd494  : out_data_ref <= 8'h44;
      11'd495  : out_data_ref <= 8'h2a;
      11'd496  : out_data_ref <= 8'he4;
      11'd497  : out_data_ref <= 8'h32;
      11'd498  : out_data_ref <= 8'h63;
      11'd499  : out_data_ref <= 8'hf9;
      11'd500  : out_data_ref <= 8'hd3;
      11'd501  : out_data_ref <= 8'h12;
      11'd502  : out_data_ref <= 8'hba;
      11'd503  : out_data_ref <= 8'hf1;
      11'd504  : out_data_ref <= 8'hd6;
      11'd505  : out_data_ref <= 8'h44;
      11'd506  : out_data_ref <= 8'h42;
      11'd507  : out_data_ref <= 8'hfd;
      11'd508  : out_data_ref <= 8'h8a;
      11'd509  : out_data_ref <= 8'hb1;
      11'd510  : out_data_ref <= 8'hf8;
      11'd511  : out_data_ref <= 8'hd7;
      11'd512  : out_data_ref <= 8'h1d;
      11'd513  : out_data_ref <= 8'h59;
      11'd514  : out_data_ref <= 8'hce;
      11'd515  : out_data_ref <= 8'h82;
      11'd516  : out_data_ref <= 8'h19;
      11'd517  : out_data_ref <= 8'h14;
      11'd518  : out_data_ref <= 8'h3e;
      11'd519  : out_data_ref <= 8'hbb;
      11'd520  : out_data_ref <= 8'hb3;
      11'd521  : out_data_ref <= 8'h8b;
      11'd522  : out_data_ref <= 8'hd9;
      11'd523  : out_data_ref <= 8'h8e;
      11'd524  : out_data_ref <= 8'h5f;
      11'd525  : out_data_ref <= 8'h37;
      11'd526  : out_data_ref <= 8'hf2;
      11'd527  : out_data_ref <= 8'h0a;
      11'd528  : out_data_ref <= 8'hb7;
      11'd529  : out_data_ref <= 8'h58;
      11'd530  : out_data_ref <= 8'h4e;
      11'd531  : out_data_ref <= 8'h82;
      11'd532  : out_data_ref <= 8'hbe;
      11'd533  : out_data_ref <= 8'ha5;
      11'd534  : out_data_ref <= 8'h13;
      11'd535  : out_data_ref <= 8'h12;
      11'd536  : out_data_ref <= 8'h31;
      11'd537  : out_data_ref <= 8'hef;
      11'd538  : out_data_ref <= 8'h6d;
      11'd539  : out_data_ref <= 8'hf8;
      11'd540  : out_data_ref <= 8'he5;
      11'd541  : out_data_ref <= 8'h11;
      11'd542  : out_data_ref <= 8'hf9;
      11'd543  : out_data_ref <= 8'ha6;
      11'd544  : out_data_ref <= 8'h2f;
      11'd545  : out_data_ref <= 8'hb4;
      11'd546  : out_data_ref <= 8'h10;
      11'd547  : out_data_ref <= 8'hfe;
      11'd548  : out_data_ref <= 8'he3;
      11'd549  : out_data_ref <= 8'h2a;
      11'd550  : out_data_ref <= 8'h16;
      11'd551  : out_data_ref <= 8'h6e;
      11'd552  : out_data_ref <= 8'hf9;
      11'd553  : out_data_ref <= 8'hef;
      11'd554  : out_data_ref <= 8'hfa;
      11'd555  : out_data_ref <= 8'h7d;
      11'd556  : out_data_ref <= 8'h30;
      11'd557  : out_data_ref <= 8'hd0;
      11'd558  : out_data_ref <= 8'hd6;
      11'd559  : out_data_ref <= 8'ha0;
      11'd560  : out_data_ref <= 8'hab;
      11'd561  : out_data_ref <= 8'hfd;
      11'd562  : out_data_ref <= 8'he3;
      11'd563  : out_data_ref <= 8'h24;
      11'd564  : out_data_ref <= 8'h87;
      11'd565  : out_data_ref <= 8'hd5;
      11'd566  : out_data_ref <= 8'heb;
      11'd567  : out_data_ref <= 8'h89;
      11'd568  : out_data_ref <= 8'hbc;
      11'd569  : out_data_ref <= 8'h54;
      11'd570  : out_data_ref <= 8'h81;
      11'd571  : out_data_ref <= 8'hef;
      11'd572  : out_data_ref <= 8'h4e;
      11'd573  : out_data_ref <= 8'he2;
      11'd574  : out_data_ref <= 8'hda;
      11'd575  : out_data_ref <= 8'h33;
      11'd576  : out_data_ref <= 8'hcb;
      11'd577  : out_data_ref <= 8'he7;
      11'd578  : out_data_ref <= 8'h32;
      11'd579  : out_data_ref <= 8'hc8;
      11'd580  : out_data_ref <= 8'h78;
      11'd581  : out_data_ref <= 8'hca;
      11'd582  : out_data_ref <= 8'hdf;
      11'd583  : out_data_ref <= 8'hc4;
      11'd584  : out_data_ref <= 8'h85;
      11'd585  : out_data_ref <= 8'h8a;
      11'd586  : out_data_ref <= 8'h0b;
      11'd587  : out_data_ref <= 8'hf4;
      11'd588  : out_data_ref <= 8'hbd;
      11'd589  : out_data_ref <= 8'h59;
      11'd590  : out_data_ref <= 8'hf2;
      11'd591  : out_data_ref <= 8'h7b;
      11'd592  : out_data_ref <= 8'h12;
      11'd593  : out_data_ref <= 8'h9c;
      11'd594  : out_data_ref <= 8'h5a;
      11'd595  : out_data_ref <= 8'hfe;
      11'd596  : out_data_ref <= 8'h60;
      11'd597  : out_data_ref <= 8'h32;
      11'd598  : out_data_ref <= 8'h7c;
      11'd599  : out_data_ref <= 8'h79;
      11'd600  : out_data_ref <= 8'h49;
      11'd601  : out_data_ref <= 8'h5a;
      11'd602  : out_data_ref <= 8'h53;
      11'd603  : out_data_ref <= 8'hf9;
      11'd604  : out_data_ref <= 8'h01;
      11'd605  : out_data_ref <= 8'hda;
      11'd606  : out_data_ref <= 8'hed;
      11'd607  : out_data_ref <= 8'hf2;
      11'd608  : out_data_ref <= 8'h71;
      11'd609  : out_data_ref <= 8'he6;
      11'd610  : out_data_ref <= 8'h40;
      11'd611  : out_data_ref <= 8'h2d;
      11'd612  : out_data_ref <= 8'h5b;
      11'd613  : out_data_ref <= 8'he7;
      11'd614  : out_data_ref <= 8'h84;
      11'd615  : out_data_ref <= 8'hf6;
      11'd616  : out_data_ref <= 8'hb3;
      11'd617  : out_data_ref <= 8'h9f;
      11'd618  : out_data_ref <= 8'hd9;
      11'd619  : out_data_ref <= 8'h88;
      11'd620  : out_data_ref <= 8'h8a;
      11'd621  : out_data_ref <= 8'h31;
      11'd622  : out_data_ref <= 8'h59;
      11'd623  : out_data_ref <= 8'h82;
      11'd624  : out_data_ref <= 8'hd9;
      11'd625  : out_data_ref <= 8'hdd;
      11'd626  : out_data_ref <= 8'h85;
      11'd627  : out_data_ref <= 8'hb0;
      11'd628  : out_data_ref <= 8'ha1;
      11'd629  : out_data_ref <= 8'h1d;
      11'd630  : out_data_ref <= 8'h43;
      11'd631  : out_data_ref <= 8'h1b;
      11'd632  : out_data_ref <= 8'hc0;
      11'd633  : out_data_ref <= 8'h8d;
      11'd634  : out_data_ref <= 8'h6e;
      11'd635  : out_data_ref <= 8'h8c;
      11'd636  : out_data_ref <= 8'h0f;
      11'd637  : out_data_ref <= 8'hac;
      11'd638  : out_data_ref <= 8'hbc;
      11'd639  : out_data_ref <= 8'h97;
      11'd640  : out_data_ref <= 8'h11;
      11'd641  : out_data_ref <= 8'he2;
      11'd642  : out_data_ref <= 8'h52;
      11'd643  : out_data_ref <= 8'h37;
      11'd644  : out_data_ref <= 8'h2d;
      11'd645  : out_data_ref <= 8'h38;
      11'd646  : out_data_ref <= 8'h6e;
      11'd647  : out_data_ref <= 8'hc4;
      11'd648  : out_data_ref <= 8'h25;
      11'd649  : out_data_ref <= 8'h39;
      11'd650  : out_data_ref <= 8'ha7;
      11'd651  : out_data_ref <= 8'h69;
      11'd652  : out_data_ref <= 8'h1f;
      11'd653  : out_data_ref <= 8'ha4;
      11'd654  : out_data_ref <= 8'hcc;
      11'd655  : out_data_ref <= 8'h40;
      11'd656  : out_data_ref <= 8'he6;
      11'd657  : out_data_ref <= 8'he4;
      11'd658  : out_data_ref <= 8'he6;
      11'd659  : out_data_ref <= 8'h4f;
      11'd660  : out_data_ref <= 8'h35;
      11'd661  : out_data_ref <= 8'h4c;
      11'd662  : out_data_ref <= 8'h12;
      11'd663  : out_data_ref <= 8'h7b;
      11'd664  : out_data_ref <= 8'hde;
      11'd665  : out_data_ref <= 8'hf2;
      11'd666  : out_data_ref <= 8'hf8;
      11'd667  : out_data_ref <= 8'h2c;
      11'd668  : out_data_ref <= 8'h45;
      11'd669  : out_data_ref <= 8'h43;
      11'd670  : out_data_ref <= 8'ha7;
      11'd671  : out_data_ref <= 8'hdf;
      11'd672  : out_data_ref <= 8'h6f;
      11'd673  : out_data_ref <= 8'h62;
      11'd674  : out_data_ref <= 8'h7e;
      11'd675  : out_data_ref <= 8'h59;
      11'd676  : out_data_ref <= 8'h71;
      11'd677  : out_data_ref <= 8'h6d;
      11'd678  : out_data_ref <= 8'hc2;
      11'd679  : out_data_ref <= 8'hcb;
      11'd680  : out_data_ref <= 8'he7;
      11'd681  : out_data_ref <= 8'had;
      11'd682  : out_data_ref <= 8'hf2;
      11'd683  : out_data_ref <= 8'hcb;
      11'd684  : out_data_ref <= 8'h24;
      11'd685  : out_data_ref <= 8'h5d;
      11'd686  : out_data_ref <= 8'hd1;
      11'd687  : out_data_ref <= 8'hcf;
      11'd688  : out_data_ref <= 8'h72;
      11'd689  : out_data_ref <= 8'h20;
      11'd690  : out_data_ref <= 8'hb6;
      11'd691  : out_data_ref <= 8'h1a;
      11'd692  : out_data_ref <= 8'h13;
      11'd693  : out_data_ref <= 8'hb0;
      11'd694  : out_data_ref <= 8'h79;
      11'd695  : out_data_ref <= 8'h61;
      11'd696  : out_data_ref <= 8'hd6;
      11'd697  : out_data_ref <= 8'h6e;
      11'd698  : out_data_ref <= 8'h21;
      11'd699  : out_data_ref <= 8'h97;
      11'd700  : out_data_ref <= 8'h98;
      11'd701  : out_data_ref <= 8'h19;
      11'd702  : out_data_ref <= 8'ha1;
      11'd703  : out_data_ref <= 8'had;
      11'd704  : out_data_ref <= 8'h61;
      11'd705  : out_data_ref <= 8'h91;
      11'd706  : out_data_ref <= 8'hf9;
      11'd707  : out_data_ref <= 8'hd3;
      11'd708  : out_data_ref <= 8'h8b;
      11'd709  : out_data_ref <= 8'hd3;
      11'd710  : out_data_ref <= 8'hf4;
      11'd711  : out_data_ref <= 8'hec;
      11'd712  : out_data_ref <= 8'hc6;
      11'd713  : out_data_ref <= 8'h31;
      11'd714  : out_data_ref <= 8'hd0;
      11'd715  : out_data_ref <= 8'hf6;
      11'd716  : out_data_ref <= 8'h61;
      11'd717  : out_data_ref <= 8'hb1;
      11'd718  : out_data_ref <= 8'h81;
      11'd719  : out_data_ref <= 8'h0b;
      11'd720  : out_data_ref <= 8'h4f;
      11'd721  : out_data_ref <= 8'ha6;
      11'd722  : out_data_ref <= 8'he4;
      11'd723  : out_data_ref <= 8'h59;
      11'd724  : out_data_ref <= 8'h34;
      11'd725  : out_data_ref <= 8'h90;
      11'd726  : out_data_ref <= 8'hdc;
      11'd727  : out_data_ref <= 8'h99;
      11'd728  : out_data_ref <= 8'h94;
      11'd729  : out_data_ref <= 8'h84;
      11'd730  : out_data_ref <= 8'hf4;
      11'd731  : out_data_ref <= 8'h73;
      11'd732  : out_data_ref <= 8'hcd;
      11'd733  : out_data_ref <= 8'h3d;
      11'd734  : out_data_ref <= 8'h64;
      11'd735  : out_data_ref <= 8'hfe;
      11'd736  : out_data_ref <= 8'hab;
      11'd737  : out_data_ref <= 8'h34;
      11'd738  : out_data_ref <= 8'hca;
      11'd739  : out_data_ref <= 8'h7b;
      11'd740  : out_data_ref <= 8'h17;
      11'd741  : out_data_ref <= 8'had;
      11'd742  : out_data_ref <= 8'ha2;
      11'd743  : out_data_ref <= 8'h19;
      11'd744  : out_data_ref <= 8'haf;
      11'd745  : out_data_ref <= 8'he7;
      11'd746  : out_data_ref <= 8'hfe;
      11'd747  : out_data_ref <= 8'h1d;
      11'd748  : out_data_ref <= 8'he5;
      11'd749  : out_data_ref <= 8'h4a;
      11'd750  : out_data_ref <= 8'had;
      11'd751  : out_data_ref <= 8'h0d;
      11'd752  : out_data_ref <= 8'h36;
      11'd753  : out_data_ref <= 8'ha8;
      11'd754  : out_data_ref <= 8'h47;
      11'd755  : out_data_ref <= 8'h59;
      11'd756  : out_data_ref <= 8'h63;
      11'd757  : out_data_ref <= 8'h6a;
      11'd758  : out_data_ref <= 8'hc3;
      11'd759  : out_data_ref <= 8'h2c;
      11'd760  : out_data_ref <= 8'hf4;
      11'd761  : out_data_ref <= 8'hbf;
      11'd762  : out_data_ref <= 8'h36;
      11'd763  : out_data_ref <= 8'hc1;
      11'd764  : out_data_ref <= 8'h7c;
      11'd765  : out_data_ref <= 8'h72;
      11'd766  : out_data_ref <= 8'haa;
      11'd767  : out_data_ref <= 8'hca;
      11'd768  : out_data_ref <= 8'h41;
      11'd769  : out_data_ref <= 8'hc0;
      11'd770  : out_data_ref <= 8'hd5;
      11'd771  : out_data_ref <= 8'h6f;
      11'd772  : out_data_ref <= 8'he2;
      11'd773  : out_data_ref <= 8'ha1;
      11'd774  : out_data_ref <= 8'h08;
      11'd775  : out_data_ref <= 8'hfc;
      11'd776  : out_data_ref <= 8'h6b;
      11'd777  : out_data_ref <= 8'hb5;
      11'd778  : out_data_ref <= 8'h43;
      11'd779  : out_data_ref <= 8'h2f;
      11'd780  : out_data_ref <= 8'h59;
      11'd781  : out_data_ref <= 8'h15;
      11'd782  : out_data_ref <= 8'h36;
      11'd783  : out_data_ref <= 8'h4c;
      11'd784  : out_data_ref <= 8'h83;
      11'd785  : out_data_ref <= 8'h0f;
      11'd786  : out_data_ref <= 8'h6a;
      11'd787  : out_data_ref <= 8'h76;
      11'd788  : out_data_ref <= 8'hd2;
      11'd789  : out_data_ref <= 8'h6a;
      11'd790  : out_data_ref <= 8'h76;
      11'd791  : out_data_ref <= 8'h88;
      11'd792  : out_data_ref <= 8'h61;
      11'd793  : out_data_ref <= 8'h51;
      11'd794  : out_data_ref <= 8'hd9;
      11'd795  : out_data_ref <= 8'h51;
      11'd796  : out_data_ref <= 8'h02;
      11'd797  : out_data_ref <= 8'h46;
      11'd798  : out_data_ref <= 8'h23;
      11'd799  : out_data_ref <= 8'he6;
      11'd800  : out_data_ref <= 8'hd7;
      11'd801  : out_data_ref <= 8'h35;
      11'd802  : out_data_ref <= 8'h6b;
      11'd803  : out_data_ref <= 8'h25;
      11'd804  : out_data_ref <= 8'hf4;
      11'd805  : out_data_ref <= 8'hd2;
      11'd806  : out_data_ref <= 8'ha2;
      11'd807  : out_data_ref <= 8'hd0;
      11'd808  : out_data_ref <= 8'h13;
      11'd809  : out_data_ref <= 8'hf9;
      11'd810  : out_data_ref <= 8'h09;
      11'd811  : out_data_ref <= 8'h28;
      11'd812  : out_data_ref <= 8'hae;
      11'd813  : out_data_ref <= 8'h3c;
      11'd814  : out_data_ref <= 8'h4b;
      11'd815  : out_data_ref <= 8'hc1;
      11'd816  : out_data_ref <= 8'hda;
      11'd817  : out_data_ref <= 8'h3e;
      11'd818  : out_data_ref <= 8'hf3;
      11'd819  : out_data_ref <= 8'hf2;
      11'd820  : out_data_ref <= 8'hd2;
      11'd821  : out_data_ref <= 8'h7d;
      11'd822  : out_data_ref <= 8'hb0;
      11'd823  : out_data_ref <= 8'ha1;
      11'd824  : out_data_ref <= 8'hff;
      11'd825  : out_data_ref <= 8'h55;
      11'd826  : out_data_ref <= 8'h90;
      11'd827  : out_data_ref <= 8'h85;
      11'd828  : out_data_ref <= 8'h6d;
      11'd829  : out_data_ref <= 8'h84;
      11'd830  : out_data_ref <= 8'h2f;
      11'd831  : out_data_ref <= 8'hfe;
      11'd832  : out_data_ref <= 8'hd5;
      11'd833  : out_data_ref <= 8'h4a;
      11'd834  : out_data_ref <= 8'h3b;
      11'd835  : out_data_ref <= 8'h9c;
      11'd836  : out_data_ref <= 8'h36;
      11'd837  : out_data_ref <= 8'hb4;
      11'd838  : out_data_ref <= 8'h10;
      11'd839  : out_data_ref <= 8'h0f;
      11'd840  : out_data_ref <= 8'hc3;
      11'd841  : out_data_ref <= 8'h38;
      11'd842  : out_data_ref <= 8'hc6;
      11'd843  : out_data_ref <= 8'h05;
      11'd844  : out_data_ref <= 8'h32;
      11'd845  : out_data_ref <= 8'had;
      11'd846  : out_data_ref <= 8'h90;
      11'd847  : out_data_ref <= 8'h4b;
      11'd848  : out_data_ref <= 8'h77;
      11'd849  : out_data_ref <= 8'h36;
      11'd850  : out_data_ref <= 8'h8d;
      11'd851  : out_data_ref <= 8'h50;
      11'd852  : out_data_ref <= 8'h6d;
      11'd853  : out_data_ref <= 8'hd4;
      11'd854  : out_data_ref <= 8'haf;
      11'd855  : out_data_ref <= 8'hba;
      11'd856  : out_data_ref <= 8'h65;
      11'd857  : out_data_ref <= 8'h0a;
      11'd858  : out_data_ref <= 8'h34;
      11'd859  : out_data_ref <= 8'hd9;
      11'd860  : out_data_ref <= 8'hc7;
      11'd861  : out_data_ref <= 8'h0e;
      11'd862  : out_data_ref <= 8'hd0;
      11'd863  : out_data_ref <= 8'haa;
      11'd864  : out_data_ref <= 8'hf1;
      11'd865  : out_data_ref <= 8'hdf;
      11'd866  : out_data_ref <= 8'h3f;
      11'd867  : out_data_ref <= 8'h4b;
      11'd868  : out_data_ref <= 8'h1b;
      11'd869  : out_data_ref <= 8'h95;
      11'd870  : out_data_ref <= 8'ha2;
      11'd871  : out_data_ref <= 8'h73;
      11'd872  : out_data_ref <= 8'h70;
      11'd873  : out_data_ref <= 8'he7;
      11'd874  : out_data_ref <= 8'h0f;
      11'd875  : out_data_ref <= 8'h4a;
      11'd876  : out_data_ref <= 8'hbf;
      11'd877  : out_data_ref <= 8'hc1;
      11'd878  : out_data_ref <= 8'h61;
      11'd879  : out_data_ref <= 8'ha6;
      11'd880  : out_data_ref <= 8'h1c;
      11'd881  : out_data_ref <= 8'h6b;
      11'd882  : out_data_ref <= 8'h25;
      11'd883  : out_data_ref <= 8'hf0;
      11'd884  : out_data_ref <= 8'hae;
      11'd885  : out_data_ref <= 8'hc8;
      11'd886  : out_data_ref <= 8'h34;
      11'd887  : out_data_ref <= 8'h9c;
      11'd888  : out_data_ref <= 8'h84;
      11'd889  : out_data_ref <= 8'h08;
      11'd890  : out_data_ref <= 8'h61;
      11'd891  : out_data_ref <= 8'hd2;
      11'd892  : out_data_ref <= 8'h9f;
      11'd893  : out_data_ref <= 8'h6e;
      11'd894  : out_data_ref <= 8'hfa;
      11'd895  : out_data_ref <= 8'h6b;
      11'd896  : out_data_ref <= 8'h9f;
      11'd897  : out_data_ref <= 8'hd1;
      11'd898  : out_data_ref <= 8'h72;
      11'd899  : out_data_ref <= 8'hf0;
      11'd900  : out_data_ref <= 8'hda;
      11'd901  : out_data_ref <= 8'h28;
      11'd902  : out_data_ref <= 8'hb9;
      11'd903  : out_data_ref <= 8'h88;
      11'd904  : out_data_ref <= 8'h87;
      11'd905  : out_data_ref <= 8'hbe;
      11'd906  : out_data_ref <= 8'h1f;
      11'd907  : out_data_ref <= 8'h6b;
      11'd908  : out_data_ref <= 8'h8a;
      11'd909  : out_data_ref <= 8'hc4;
      11'd910  : out_data_ref <= 8'h95;
      11'd911  : out_data_ref <= 8'hfd;
      11'd912  : out_data_ref <= 8'h6a;
      11'd913  : out_data_ref <= 8'h54;
      11'd914  : out_data_ref <= 8'h47;
      11'd915  : out_data_ref <= 8'hdc;
      11'd916  : out_data_ref <= 8'h9a;
      11'd917  : out_data_ref <= 8'h0d;
      11'd918  : out_data_ref <= 8'h57;
      11'd919  : out_data_ref <= 8'h9c;
      11'd920  : out_data_ref <= 8'hc8;
      11'd921  : out_data_ref <= 8'h9f;
      11'd922  : out_data_ref <= 8'h37;
      11'd923  : out_data_ref <= 8'h9d;
      11'd924  : out_data_ref <= 8'h4c;
      11'd925  : out_data_ref <= 8'ha6;
      11'd926  : out_data_ref <= 8'h87;
      11'd927  : out_data_ref <= 8'he6;
      11'd928  : out_data_ref <= 8'h1c;
      11'd929  : out_data_ref <= 8'h67;
      11'd930  : out_data_ref <= 8'h87;
      11'd931  : out_data_ref <= 8'h68;
      11'd932  : out_data_ref <= 8'h98;
      11'd933  : out_data_ref <= 8'hec;
      11'd934  : out_data_ref <= 8'h2d;
      11'd935  : out_data_ref <= 8'h45;
      11'd936  : out_data_ref <= 8'hdf;
      11'd937  : out_data_ref <= 8'h4a;
      11'd938  : out_data_ref <= 8'hb3;
      11'd939  : out_data_ref <= 8'h75;
      11'd940  : out_data_ref <= 8'he1;
      11'd941  : out_data_ref <= 8'h6b;
      11'd942  : out_data_ref <= 8'h1d;
      11'd943  : out_data_ref <= 8'hd6;
      11'd944  : out_data_ref <= 8'hfc;
      11'd945  : out_data_ref <= 8'h6e;
      11'd946  : out_data_ref <= 8'h3f;
      11'd947  : out_data_ref <= 8'h8e;
      11'd948  : out_data_ref <= 8'h72;
      11'd949  : out_data_ref <= 8'h0c;
      11'd950  : out_data_ref <= 8'h45;
      11'd951  : out_data_ref <= 8'hf8;
      11'd952  : out_data_ref <= 8'ha6;
      11'd953  : out_data_ref <= 8'h35;
      11'd954  : out_data_ref <= 8'h8a;
      11'd955  : out_data_ref <= 8'h7a;
      11'd956  : out_data_ref <= 8'h21;
      11'd957  : out_data_ref <= 8'h1c;
      11'd958  : out_data_ref <= 8'h52;
      11'd959  : out_data_ref <= 8'hc6;
      11'd960  : out_data_ref <= 8'h8c;
      11'd961  : out_data_ref <= 8'h9d;
      11'd962  : out_data_ref <= 8'he4;
      11'd963  : out_data_ref <= 8'h07;
      11'd964  : out_data_ref <= 8'hb9;
      11'd965  : out_data_ref <= 8'h8e;
      11'd966  : out_data_ref <= 8'h74;
      11'd967  : out_data_ref <= 8'h3e;
      11'd968  : out_data_ref <= 8'h46;
      11'd969  : out_data_ref <= 8'h97;
      11'd970  : out_data_ref <= 8'h30;
      11'd971  : out_data_ref <= 8'h6f;
      11'd972  : out_data_ref <= 8'hc4;
      11'd973  : out_data_ref <= 8'h3f;
      11'd974  : out_data_ref <= 8'h7a;
      11'd975  : out_data_ref <= 8'h9f;
      11'd976  : out_data_ref <= 8'ha6;
      11'd977  : out_data_ref <= 8'h6c;
      11'd978  : out_data_ref <= 8'h41;
      11'd979  : out_data_ref <= 8'hb8;
      11'd980  : out_data_ref <= 8'hdf;
      11'd981  : out_data_ref <= 8'ha8;
      11'd982  : out_data_ref <= 8'h6f;
      11'd983  : out_data_ref <= 8'he6;
      11'd984  : out_data_ref <= 8'ha6;
      11'd985  : out_data_ref <= 8'he5;
      11'd986  : out_data_ref <= 8'h0c;
      11'd987  : out_data_ref <= 8'h52;
      11'd988  : out_data_ref <= 8'hd9;
      11'd989  : out_data_ref <= 8'h46;
      11'd990  : out_data_ref <= 8'h35;
      11'd991  : out_data_ref <= 8'h9e;
      11'd992  : out_data_ref <= 8'h7d;
      11'd993  : out_data_ref <= 8'he5;
      11'd994  : out_data_ref <= 8'h14;
      11'd995  : out_data_ref <= 8'h2f;
      11'd996  : out_data_ref <= 8'he5;
      11'd997  : out_data_ref <= 8'h3e;
      11'd998  : out_data_ref <= 8'h3d;
      11'd999  : out_data_ref <= 8'hee;
      11'd1000 : out_data_ref <= 8'h32;
      11'd1001 : out_data_ref <= 8'h18;
      11'd1002 : out_data_ref <= 8'h8f;
      11'd1003 : out_data_ref <= 8'h11;
      11'd1004 : out_data_ref <= 8'ha9;
      11'd1005 : out_data_ref <= 8'ha5;
      11'd1006 : out_data_ref <= 8'he7;
      11'd1007 : out_data_ref <= 8'h87;
      11'd1008 : out_data_ref <= 8'hcb;
      11'd1009 : out_data_ref <= 8'h3a;
      11'd1010 : out_data_ref <= 8'h20;
      11'd1011 : out_data_ref <= 8'hd2;
      11'd1012 : out_data_ref <= 8'h61;
      11'd1013 : out_data_ref <= 8'h38;
      11'd1014 : out_data_ref <= 8'hd6;
      11'd1015 : out_data_ref <= 8'hfd;
      11'd1016 : out_data_ref <= 8'h15;
      11'd1017 : out_data_ref <= 8'he1;
      11'd1018 : out_data_ref <= 8'h4a;
      11'd1019 : out_data_ref <= 8'h73;
      11'd1020 : out_data_ref <= 8'hda;
      11'd1021 : out_data_ref <= 8'h5a;
      11'd1022 : out_data_ref <= 8'ha9;
      11'd1023 : out_data_ref <= 8'h05;
      11'd1024 : out_data_ref <= 8'hfd;
      11'd1025 : out_data_ref <= 8'h66;
      11'd1026 : out_data_ref <= 8'h50;
      11'd1027 : out_data_ref <= 8'h40;
      11'd1028 : out_data_ref <= 8'hcc;
      11'd1029 : out_data_ref <= 8'h93;
      11'd1030 : out_data_ref <= 8'h9c;
      11'd1031 : out_data_ref <= 8'h2d;
      11'd1032 : out_data_ref <= 8'ha6;
      11'd1033 : out_data_ref <= 8'h83;
      11'd1034 : out_data_ref <= 8'h6f;
      11'd1035 : out_data_ref <= 8'h04;
      11'd1036 : out_data_ref <= 8'hed;
      11'd1037 : out_data_ref <= 8'h8b;
      11'd1038 : out_data_ref <= 8'h8c;
      11'd1039 : out_data_ref <= 8'h9f;
      11'd1040 : out_data_ref <= 8'h27;
      11'd1041 : out_data_ref <= 8'h72;
      11'd1042 : out_data_ref <= 8'h09;
      11'd1043 : out_data_ref <= 8'h20;
      11'd1044 : out_data_ref <= 8'h10;
      11'd1045 : out_data_ref <= 8'hfc;
      11'd1046 : out_data_ref <= 8'h92;
      11'd1047 : out_data_ref <= 8'hbd;
      11'd1048 : out_data_ref <= 8'h35;
      11'd1049 : out_data_ref <= 8'hdd;
      11'd1050 : out_data_ref <= 8'h40;
      11'd1051 : out_data_ref <= 8'h8c;
      11'd1052 : out_data_ref <= 8'h55;
      11'd1053 : out_data_ref <= 8'h43;
      11'd1054 : out_data_ref <= 8'hc5;
      11'd1055 : out_data_ref <= 8'hfb;
      11'd1056 : out_data_ref <= 8'h8d;
      11'd1057 : out_data_ref <= 8'hd8;
      11'd1058 : out_data_ref <= 8'hf4;
      11'd1059 : out_data_ref <= 8'h43;
      11'd1060 : out_data_ref <= 8'h4c;
      11'd1061 : out_data_ref <= 8'hf1;
      11'd1062 : out_data_ref <= 8'h1b;
      11'd1063 : out_data_ref <= 8'hd2;
      11'd1064 : out_data_ref <= 8'h8a;
      11'd1065 : out_data_ref <= 8'hb2;
      11'd1066 : out_data_ref <= 8'hb4;
      11'd1067 : out_data_ref <= 8'h65;
      11'd1068 : out_data_ref <= 8'h49;
      11'd1069 : out_data_ref <= 8'hbb;
      11'd1070 : out_data_ref <= 8'h53;
      11'd1071 : out_data_ref <= 8'hfa;
      11'd1072 : out_data_ref <= 8'h59;
      11'd1073 : out_data_ref <= 8'h52;
      11'd1074 : out_data_ref <= 8'hc6;
      11'd1075 : out_data_ref <= 8'hfd;
      11'd1076 : out_data_ref <= 8'hd7;
      11'd1077 : out_data_ref <= 8'h7c;
      11'd1078 : out_data_ref <= 8'h44;
      11'd1079 : out_data_ref <= 8'h07;
      11'd1080 : out_data_ref <= 8'he5;
      11'd1081 : out_data_ref <= 8'h9d;
      11'd1082 : out_data_ref <= 8'h10;
      11'd1083 : out_data_ref <= 8'ha6;
      11'd1084 : out_data_ref <= 8'he7;
      11'd1085 : out_data_ref <= 8'hf2;
      11'd1086 : out_data_ref <= 8'h57;
      11'd1087 : out_data_ref <= 8'h7a;
      11'd1088 : out_data_ref <= 8'hb5;
      11'd1089 : out_data_ref <= 8'h41;
      11'd1090 : out_data_ref <= 8'hc5;
      11'd1091 : out_data_ref <= 8'h9e;
      11'd1092 : out_data_ref <= 8'hb6;
      11'd1093 : out_data_ref <= 8'hc9;
      11'd1094 : out_data_ref <= 8'h14;
      11'd1095 : out_data_ref <= 8'h3f;
      11'd1096 : out_data_ref <= 8'h5d;
      11'd1097 : out_data_ref <= 8'hcd;
      11'd1098 : out_data_ref <= 8'h5f;
      11'd1099 : out_data_ref <= 8'h10;
      11'd1100 : out_data_ref <= 8'h24;
      11'd1101 : out_data_ref <= 8'h71;
      11'd1102 : out_data_ref <= 8'hea;
      11'd1103 : out_data_ref <= 8'h70;
      11'd1104 : out_data_ref <= 8'h10;
      11'd1105 : out_data_ref <= 8'hc8;
      11'd1106 : out_data_ref <= 8'hf2;
      11'd1107 : out_data_ref <= 8'h32;
      11'd1108 : out_data_ref <= 8'h64;
      11'd1109 : out_data_ref <= 8'h3f;
      11'd1110 : out_data_ref <= 8'h11;
      11'd1111 : out_data_ref <= 8'hba;
      11'd1112 : out_data_ref <= 8'he3;
      11'd1113 : out_data_ref <= 8'h1c;
      11'd1114 : out_data_ref <= 8'hbb;
      11'd1115 : out_data_ref <= 8'h9e;
      11'd1116 : out_data_ref <= 8'hb9;
      11'd1117 : out_data_ref <= 8'he0;
      11'd1118 : out_data_ref <= 8'hb2;
      11'd1119 : out_data_ref <= 8'hc5;
      11'd1120 : out_data_ref <= 8'hfa;
      11'd1121 : out_data_ref <= 8'h2c;
      11'd1122 : out_data_ref <= 8'h5a;
      11'd1123 : out_data_ref <= 8'h78;
      11'd1124 : out_data_ref <= 8'h8a;
      11'd1125 : out_data_ref <= 8'h68;
      11'd1126 : out_data_ref <= 8'h0b;
      11'd1127 : out_data_ref <= 8'hf1;
      11'd1128 : out_data_ref <= 8'h5e;
      11'd1129 : out_data_ref <= 8'h56;
      11'd1130 : out_data_ref <= 8'h8c;
      11'd1131 : out_data_ref <= 8'h42;
      11'd1132 : out_data_ref <= 8'h5a;
      11'd1133 : out_data_ref <= 8'h39;
      11'd1134 : out_data_ref <= 8'h55;
      11'd1135 : out_data_ref <= 8'hc5;
      11'd1136 : out_data_ref <= 8'h72;
      11'd1137 : out_data_ref <= 8'h40;
      11'd1138 : out_data_ref <= 8'h27;
      11'd1139 : out_data_ref <= 8'he5;
      11'd1140 : out_data_ref <= 8'h21;
      11'd1141 : out_data_ref <= 8'h12;
      11'd1142 : out_data_ref <= 8'h7b;
      11'd1143 : out_data_ref <= 8'h1d;
      11'd1144 : out_data_ref <= 8'h4b;
      11'd1145 : out_data_ref <= 8'hac;
      11'd1146 : out_data_ref <= 8'h12;
      11'd1147 : out_data_ref <= 8'h71;
      11'd1148 : out_data_ref <= 8'h82;
      11'd1149 : out_data_ref <= 8'hc7;
      11'd1150 : out_data_ref <= 8'h16;
      11'd1151 : out_data_ref <= 8'h97;
      11'd1152 : out_data_ref <= 8'h61;
      11'd1153 : out_data_ref <= 8'h02;
      11'd1154 : out_data_ref <= 8'hd0;
      11'd1155 : out_data_ref <= 8'hdd;
      11'd1156 : out_data_ref <= 8'he8;
      11'd1157 : out_data_ref <= 8'h16;
      11'd1158 : out_data_ref <= 8'hab;
      11'd1159 : out_data_ref <= 8'h4e;
      11'd1160 : out_data_ref <= 8'h8e;
      11'd1161 : out_data_ref <= 8'h3f;
      11'd1162 : out_data_ref <= 8'he4;
      11'd1163 : out_data_ref <= 8'h8e;
      11'd1164 : out_data_ref <= 8'hb9;
      11'd1165 : out_data_ref <= 8'h28;
      11'd1166 : out_data_ref <= 8'h9b;
      11'd1167 : out_data_ref <= 8'hbf;
      11'd1168 : out_data_ref <= 8'h47;
      11'd1169 : out_data_ref <= 8'h79;
      11'd1170 : out_data_ref <= 8'h17;
      11'd1171 : out_data_ref <= 8'hbe;
      11'd1172 : out_data_ref <= 8'h58;
      11'd1173 : out_data_ref <= 8'h04;
      11'd1174 : out_data_ref <= 8'h4e;
      11'd1175 : out_data_ref <= 8'h97;
      11'd1176 : out_data_ref <= 8'hc7;
      11'd1177 : out_data_ref <= 8'h0d;
      11'd1178 : out_data_ref <= 8'haf;
      11'd1179 : out_data_ref <= 8'hbe;
      11'd1180 : out_data_ref <= 8'he9;
      11'd1181 : out_data_ref <= 8'ha3;
      11'd1182 : out_data_ref <= 8'h77;
      11'd1183 : out_data_ref <= 8'h80;
      11'd1184 : out_data_ref <= 8'hcf;
      11'd1185 : out_data_ref <= 8'h94;
      11'd1186 : out_data_ref <= 8'hc9;
      11'd1187 : out_data_ref <= 8'hd8;
      11'd1188 : out_data_ref <= 8'h30;
      11'd1189 : out_data_ref <= 8'h89;
      11'd1190 : out_data_ref <= 8'h0a;
      11'd1191 : out_data_ref <= 8'h33;
      11'd1192 : out_data_ref <= 8'hc1;
      11'd1193 : out_data_ref <= 8'h12;
      11'd1194 : out_data_ref <= 8'h50;
      11'd1195 : out_data_ref <= 8'h14;
      11'd1196 : out_data_ref <= 8'hf2;
      11'd1197 : out_data_ref <= 8'hf9;
      11'd1198 : out_data_ref <= 8'hda;
      11'd1199 : out_data_ref <= 8'h87;
      11'd1200 : out_data_ref <= 8'hdf;
      11'd1201 : out_data_ref <= 8'h36;
      11'd1202 : out_data_ref <= 8'hcb;
      11'd1203 : out_data_ref <= 8'h26;
      11'd1204 : out_data_ref <= 8'h7a;
      11'd1205 : out_data_ref <= 8'h33;
      11'd1206 : out_data_ref <= 8'h8d;
      11'd1207 : out_data_ref <= 8'h66;
      11'd1208 : out_data_ref <= 8'hf2;
      11'd1209 : out_data_ref <= 8'h9c;
      11'd1210 : out_data_ref <= 8'he2;
      11'd1211 : out_data_ref <= 8'h89;
      11'd1212 : out_data_ref <= 8'h3a;
      11'd1213 : out_data_ref <= 8'h11;
      11'd1214 : out_data_ref <= 8'h74;
      11'd1215 : out_data_ref <= 8'h5d;
      11'd1216 : out_data_ref <= 8'ha1;
      11'd1217 : out_data_ref <= 8'h08;
      11'd1218 : out_data_ref <= 8'hb9;
      11'd1219 : out_data_ref <= 8'hf0;
      11'd1220 : out_data_ref <= 8'h5e;
      11'd1221 : out_data_ref <= 8'h40;
      11'd1222 : out_data_ref <= 8'hca;
      11'd1223 : out_data_ref <= 8'h46;
      11'd1224 : out_data_ref <= 8'hd9;
      11'd1225 : out_data_ref <= 8'h65;
      11'd1226 : out_data_ref <= 8'hed;
      11'd1227 : out_data_ref <= 8'h7a;
      11'd1228 : out_data_ref <= 8'h18;
      11'd1229 : out_data_ref <= 8'h26;
      11'd1230 : out_data_ref <= 8'h9b;
      11'd1231 : out_data_ref <= 8'h56;
      11'd1232 : out_data_ref <= 8'hf3;
      11'd1233 : out_data_ref <= 8'h7d;
      11'd1234 : out_data_ref <= 8'hcb;
      11'd1235 : out_data_ref <= 8'h2a;
      11'd1236 : out_data_ref <= 8'h96;
      11'd1237 : out_data_ref <= 8'h37;
      11'd1238 : out_data_ref <= 8'ha8;
      11'd1239 : out_data_ref <= 8'hb9;
      11'd1240 : out_data_ref <= 8'h69;
      11'd1241 : out_data_ref <= 8'h24;
      11'd1242 : out_data_ref <= 8'hcd;
      11'd1243 : out_data_ref <= 8'h29;
      11'd1244 : out_data_ref <= 8'hb9;
      11'd1245 : out_data_ref <= 8'h70;
      11'd1246 : out_data_ref <= 8'h8c;
      11'd1247 : out_data_ref <= 8'h50;
      11'd1248 : out_data_ref <= 8'hcc;
      11'd1249 : out_data_ref <= 8'h14;
      11'd1250 : out_data_ref <= 8'hab;
      11'd1251 : out_data_ref <= 8'hbd;
      11'd1252 : out_data_ref <= 8'h2c;
      11'd1253 : out_data_ref <= 8'hb4;
      11'd1254 : out_data_ref <= 8'hca;
      11'd1255 : out_data_ref <= 8'h0d;
      11'd1256 : out_data_ref <= 8'h9d;
      11'd1257 : out_data_ref <= 8'h26;
      11'd1258 : out_data_ref <= 8'h4d;
      11'd1259 : out_data_ref <= 8'h0c;
      11'd1260 : out_data_ref <= 8'h3d;
      11'd1261 : out_data_ref <= 8'haa;
      11'd1262 : out_data_ref <= 8'hf0;
      11'd1263 : out_data_ref <= 8'h8e;
      11'd1264 : out_data_ref <= 8'h16;
      11'd1265 : out_data_ref <= 8'h9e;
      11'd1266 : out_data_ref <= 8'h83;
      11'd1267 : out_data_ref <= 8'hd8;
      11'd1268 : out_data_ref <= 8'hff;
      11'd1269 : out_data_ref <= 8'hdb;
      11'd1270 : out_data_ref <= 8'h11;
      11'd1271 : out_data_ref <= 8'h5f;
      11'd1272 : out_data_ref <= 8'h83;
      11'd1273 : out_data_ref <= 8'h92;
      11'd1274 : out_data_ref <= 8'hfd;
      11'd1275 : out_data_ref <= 8'h32;
      11'd1276 : out_data_ref <= 8'h65;
      11'd1277 : out_data_ref <= 8'h98;
      11'd1278 : out_data_ref <= 8'h4d;
      11'd1279 : out_data_ref <= 8'h23;
      11'd1280 : out_data_ref <= 8'h80;
      11'd1281 : out_data_ref <= 8'hb3;
      11'd1282 : out_data_ref <= 8'h59;
      11'd1283 : out_data_ref <= 8'h89;
      11'd1284 : out_data_ref <= 8'h55;
      11'd1285 : out_data_ref <= 8'ha7;
      11'd1286 : out_data_ref <= 8'hb3;
      11'd1287 : out_data_ref <= 8'hb2;
      11'd1288 : out_data_ref <= 8'h8b;
      11'd1289 : out_data_ref <= 8'hf2;
      11'd1290 : out_data_ref <= 8'hdd;
      11'd1291 : out_data_ref <= 8'h06;
      11'd1292 : out_data_ref <= 8'h92;
      11'd1293 : out_data_ref <= 8'h0a;
      11'd1294 : out_data_ref <= 8'h2f;
      11'd1295 : out_data_ref <= 8'hf0;
      11'd1296 : out_data_ref <= 8'hdd;
      11'd1297 : out_data_ref <= 8'hb7;
      11'd1298 : out_data_ref <= 8'hef;
      11'd1299 : out_data_ref <= 8'h96;
      11'd1300 : out_data_ref <= 8'hf1;
      11'd1301 : out_data_ref <= 8'h70;
      11'd1302 : out_data_ref <= 8'haf;
      11'd1303 : out_data_ref <= 8'h03;
      11'd1304 : out_data_ref <= 8'hd1;
      11'd1305 : out_data_ref <= 8'h9f;
      11'd1306 : out_data_ref <= 8'ha2;
      11'd1307 : out_data_ref <= 8'hca;
      11'd1308 : out_data_ref <= 8'hbe;
      11'd1309 : out_data_ref <= 8'ha2;
      11'd1310 : out_data_ref <= 8'h3a;
      11'd1311 : out_data_ref <= 8'ha3;
      11'd1312 : out_data_ref <= 8'hce;
      11'd1313 : out_data_ref <= 8'h97;
      11'd1314 : out_data_ref <= 8'h5d;
      11'd1315 : out_data_ref <= 8'he4;
      11'd1316 : out_data_ref <= 8'hcc;
      11'd1317 : out_data_ref <= 8'h01;
      11'd1318 : out_data_ref <= 8'he3;
      11'd1319 : out_data_ref <= 8'h7d;
      11'd1320 : out_data_ref <= 8'h17;
      11'd1321 : out_data_ref <= 8'he8;
      11'd1322 : out_data_ref <= 8'he3;
      11'd1323 : out_data_ref <= 8'hec;
      11'd1324 : out_data_ref <= 8'h13;
      11'd1325 : out_data_ref <= 8'h01;
      11'd1326 : out_data_ref <= 8'h86;
      11'd1327 : out_data_ref <= 8'h3a;
      11'd1328 : out_data_ref <= 8'h6a;
      11'd1329 : out_data_ref <= 8'h4e;
      11'd1330 : out_data_ref <= 8'h24;
      11'd1331 : out_data_ref <= 8'h18;
      11'd1332 : out_data_ref <= 8'h8f;
      11'd1333 : out_data_ref <= 8'h17;
      11'd1334 : out_data_ref <= 8'h65;
      11'd1335 : out_data_ref <= 8'haa;
      11'd1336 : out_data_ref <= 8'hfa;
      11'd1337 : out_data_ref <= 8'h75;
      11'd1338 : out_data_ref <= 8'hf9;
      11'd1339 : out_data_ref <= 8'hdd;
      11'd1340 : out_data_ref <= 8'hdd;
      11'd1341 : out_data_ref <= 8'h64;
      11'd1342 : out_data_ref <= 8'hd3;
      11'd1343 : out_data_ref <= 8'haf;
      11'd1344 : out_data_ref <= 8'he7;
      11'd1345 : out_data_ref <= 8'h19;
      11'd1346 : out_data_ref <= 8'h90;
      11'd1347 : out_data_ref <= 8'hb1;
      11'd1348 : out_data_ref <= 8'hdc;
      11'd1349 : out_data_ref <= 8'h4a;
      11'd1350 : out_data_ref <= 8'h6a;
      11'd1351 : out_data_ref <= 8'h05;
      11'd1352 : out_data_ref <= 8'h7e;
      11'd1353 : out_data_ref <= 8'h56;
      11'd1354 : out_data_ref <= 8'h33;
      11'd1355 : out_data_ref <= 8'he1;
      11'd1356 : out_data_ref <= 8'hf4;
      11'd1357 : out_data_ref <= 8'h40;
      11'd1358 : out_data_ref <= 8'h97;
      11'd1359 : out_data_ref <= 8'hc1;
      11'd1360 : out_data_ref <= 8'hb7;
      11'd1361 : out_data_ref <= 8'hd9;
      11'd1362 : out_data_ref <= 8'h94;
      11'd1363 : out_data_ref <= 8'h3a;
      11'd1364 : out_data_ref <= 8'h3c;
      11'd1365 : out_data_ref <= 8'h79;
      11'd1366 : out_data_ref <= 8'h79;
      11'd1367 : out_data_ref <= 8'ha7;
      11'd1368 : out_data_ref <= 8'h96;
      11'd1369 : out_data_ref <= 8'hdb;
      11'd1370 : out_data_ref <= 8'h67;
      11'd1371 : out_data_ref <= 8'h6d;
      11'd1372 : out_data_ref <= 8'ha3;
      11'd1373 : out_data_ref <= 8'h4e;
      11'd1374 : out_data_ref <= 8'h6b;
      11'd1375 : out_data_ref <= 8'hd6;
      11'd1376 : out_data_ref <= 8'h88;
      11'd1377 : out_data_ref <= 8'h3c;
      11'd1378 : out_data_ref <= 8'h43;
      11'd1379 : out_data_ref <= 8'hc0;
      11'd1380 : out_data_ref <= 8'h43;
      11'd1381 : out_data_ref <= 8'h43;
      11'd1382 : out_data_ref <= 8'h57;
      11'd1383 : out_data_ref <= 8'hee;
      11'd1384 : out_data_ref <= 8'hc0;
      11'd1385 : out_data_ref <= 8'hf7;
      11'd1386 : out_data_ref <= 8'h53;
      11'd1387 : out_data_ref <= 8'h00;
      11'd1388 : out_data_ref <= 8'h1f;
      11'd1389 : out_data_ref <= 8'hc1;
      11'd1390 : out_data_ref <= 8'haf;
      11'd1391 : out_data_ref <= 8'h4f;
      11'd1392 : out_data_ref <= 8'he4;
      11'd1393 : out_data_ref <= 8'he4;
      11'd1394 : out_data_ref <= 8'hf5;
      11'd1395 : out_data_ref <= 8'h94;
      11'd1396 : out_data_ref <= 8'hf6;
      11'd1397 : out_data_ref <= 8'haf;
      11'd1398 : out_data_ref <= 8'hcc;
      11'd1399 : out_data_ref <= 8'h81;
      11'd1400 : out_data_ref <= 8'h32;
      11'd1401 : out_data_ref <= 8'hc4;
      11'd1402 : out_data_ref <= 8'h4b;
      11'd1403 : out_data_ref <= 8'hdd;
      11'd1404 : out_data_ref <= 8'h95;
      11'd1405 : out_data_ref <= 8'ha1;
      11'd1406 : out_data_ref <= 8'hfa;
      11'd1407 : out_data_ref <= 8'h7d;
      11'd1408 : out_data_ref <= 8'h2e;
      11'd1409 : out_data_ref <= 8'hef;
      11'd1410 : out_data_ref <= 8'h0e;
      11'd1411 : out_data_ref <= 8'h71;
      11'd1412 : out_data_ref <= 8'hb4;
      11'd1413 : out_data_ref <= 8'h6c;
      11'd1414 : out_data_ref <= 8'h3c;
      11'd1415 : out_data_ref <= 8'h23;
      11'd1416 : out_data_ref <= 8'h8d;
      11'd1417 : out_data_ref <= 8'h88;
      11'd1418 : out_data_ref <= 8'h94;
      11'd1419 : out_data_ref <= 8'h96;
      11'd1420 : out_data_ref <= 8'h39;
      11'd1421 : out_data_ref <= 8'h6a;
      11'd1422 : out_data_ref <= 8'h8f;
      11'd1423 : out_data_ref <= 8'h5f;
      11'd1424 : out_data_ref <= 8'h42;
      11'd1425 : out_data_ref <= 8'hc1;
      11'd1426 : out_data_ref <= 8'h94;
      11'd1427 : out_data_ref <= 8'hd9;
      11'd1428 : out_data_ref <= 8'hb3;
      11'd1429 : out_data_ref <= 8'h33;
      11'd1430 : out_data_ref <= 8'hf2;
      11'd1431 : out_data_ref <= 8'h49;
      11'd1432 : out_data_ref <= 8'h10;
      11'd1433 : out_data_ref <= 8'h53;
      11'd1434 : out_data_ref <= 8'h8a;
      11'd1435 : out_data_ref <= 8'hf8;
      11'd1436 : out_data_ref <= 8'h43;
      11'd1437 : out_data_ref <= 8'hc9;
      11'd1438 : out_data_ref <= 8'h3e;
      11'd1439 : out_data_ref <= 8'h79;
      11'd1440 : out_data_ref <= 8'h2e;
      11'd1441 : out_data_ref <= 8'h10;
      11'd1442 : out_data_ref <= 8'hfc;
      11'd1443 : out_data_ref <= 8'hd2;
      11'd1444 : out_data_ref <= 8'h50;
      11'd1445 : out_data_ref <= 8'hd5;
      11'd1446 : out_data_ref <= 8'ha8;
      11'd1447 : out_data_ref <= 8'h21;
      11'd1448 : out_data_ref <= 8'hdc;
      11'd1449 : out_data_ref <= 8'h70;
      11'd1450 : out_data_ref <= 8'h2c;
      11'd1451 : out_data_ref <= 8'hae;
      11'd1452 : out_data_ref <= 8'h00;
      11'd1453 : out_data_ref <= 8'h7a;
      11'd1454 : out_data_ref <= 8'h6b;
      11'd1455 : out_data_ref <= 8'hcd;
      11'd1456 : out_data_ref <= 8'hcc;
      11'd1457 : out_data_ref <= 8'hfb;
      11'd1458 : out_data_ref <= 8'h34;
      11'd1459 : out_data_ref <= 8'h78;
      11'd1460 : out_data_ref <= 8'h8f;
      11'd1461 : out_data_ref <= 8'h8a;
      11'd1462 : out_data_ref <= 8'h1a;
      11'd1463 : out_data_ref <= 8'h7e;
      11'd1464 : out_data_ref <= 8'h9c;
      11'd1465 : out_data_ref <= 8'h26;
      11'd1466 : out_data_ref <= 8'h19;
      11'd1467 : out_data_ref <= 8'h71;
      11'd1468 : out_data_ref <= 8'h38;
      11'd1469 : out_data_ref <= 8'h1f;
      11'd1470 : out_data_ref <= 8'h60;
      11'd1471 : out_data_ref <= 8'h56;
      11'd1472 : out_data_ref <= 8'hde;
      11'd1473 : out_data_ref <= 8'h61;
      11'd1474 : out_data_ref <= 8'h89;
      11'd1475 : out_data_ref <= 8'hd3;
      11'd1476 : out_data_ref <= 8'hc0;
      11'd1477 : out_data_ref <= 8'h6b;
      11'd1478 : out_data_ref <= 8'h3d;
      11'd1479 : out_data_ref <= 8'hf0;
      11'd1480 : out_data_ref <= 8'h1f;
      11'd1481 : out_data_ref <= 8'h5a;
      11'd1482 : out_data_ref <= 8'h0a;
      11'd1483 : out_data_ref <= 8'hd1;
      11'd1484 : out_data_ref <= 8'hdb;
      11'd1485 : out_data_ref <= 8'ha5;
      11'd1486 : out_data_ref <= 8'h24;
      11'd1487 : out_data_ref <= 8'h66;
      11'd1488 : out_data_ref <= 8'hc0;
      11'd1489 : out_data_ref <= 8'h4f;
      11'd1490 : out_data_ref <= 8'h61;
      11'd1491 : out_data_ref <= 8'h5e;
      11'd1492 : out_data_ref <= 8'h2b;
      11'd1493 : out_data_ref <= 8'h45;
      11'd1494 : out_data_ref <= 8'hc4;
      11'd1495 : out_data_ref <= 8'hc1;
      11'd1496 : out_data_ref <= 8'h1f;
      11'd1497 : out_data_ref <= 8'he1;
      11'd1498 : out_data_ref <= 8'h3c;
      11'd1499 : out_data_ref <= 8'ha0;
      11'd1500 : out_data_ref <= 8'had;
      11'd1501 : out_data_ref <= 8'h74;
      11'd1502 : out_data_ref <= 8'hf7;
      11'd1503 : out_data_ref <= 8'h9c;
      11'd1504 : out_data_ref <= 8'h18;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
