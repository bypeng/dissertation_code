module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd857;
  localparam R_DEPTH = 'd10;
  localparam B_LEN = 'd1322;
  localparam B_DEPTH = 'd11;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [13: 0] in_data;
  input      [10: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 14'h0e8b; // 'd3723
      10'd1    : in_data <= 14'h0ce7; // 'd3303
      10'd2    : in_data <= 14'h0fd1; // 'd4049
      10'd3    : in_data <= 14'h07f1; // 'd2033
      10'd4    : in_data <= 14'h0df7; // 'd3575
      10'd5    : in_data <= 14'h08df; // 'd2271
      10'd6    : in_data <= 14'h0bcd; // 'd3021
      10'd7    : in_data <= 14'h0285; // 'd645
      10'd8    : in_data <= 14'h0cdc; // 'd3292
      10'd9    : in_data <= 14'h0424; // 'd1060
      10'd10   : in_data <= 14'h0f73; // 'd3955
      10'd11   : in_data <= 14'h0d04; // 'd3332
      10'd12   : in_data <= 14'h0fee; // 'd4078
      10'd13   : in_data <= 14'h00a5; // 'd165
      10'd14   : in_data <= 14'h00bd; // 'd189
      10'd15   : in_data <= 14'h0858; // 'd2136
      10'd16   : in_data <= 14'h123b; // 'd4667
      10'd17   : in_data <= 14'h03a6; // 'd934
      10'd18   : in_data <= 14'h11e0; // 'd4576
      10'd19   : in_data <= 14'h0a0b; // 'd2571
      10'd20   : in_data <= 14'h1187; // 'd4487
      10'd21   : in_data <= 14'h13e6; // 'd5094
      10'd22   : in_data <= 14'h0552; // 'd1362
      10'd23   : in_data <= 14'h0993; // 'd2451
      10'd24   : in_data <= 14'h0b01; // 'd2817
      10'd25   : in_data <= 14'h095b; // 'd2395
      10'd26   : in_data <= 14'h0342; // 'd834
      10'd27   : in_data <= 14'h0e4a; // 'd3658
      10'd28   : in_data <= 14'h026c; // 'd620
      10'd29   : in_data <= 14'h05bb; // 'd1467
      10'd30   : in_data <= 14'h123e; // 'd4670
      10'd31   : in_data <= 14'h074a; // 'd1866
      10'd32   : in_data <= 14'h0607; // 'd1543
      10'd33   : in_data <= 14'h04c0; // 'd1216
      10'd34   : in_data <= 14'h121d; // 'd4637
      10'd35   : in_data <= 14'h0848; // 'd2120
      10'd36   : in_data <= 14'h001e; // 'd30
      10'd37   : in_data <= 14'h0cdf; // 'd3295
      10'd38   : in_data <= 14'h0879; // 'd2169
      10'd39   : in_data <= 14'h1282; // 'd4738
      10'd40   : in_data <= 14'h1244; // 'd4676
      10'd41   : in_data <= 14'h13b6; // 'd5046
      10'd42   : in_data <= 14'h0abe; // 'd2750
      10'd43   : in_data <= 14'h0b3c; // 'd2876
      10'd44   : in_data <= 14'h0ff8; // 'd4088
      10'd45   : in_data <= 14'h0565; // 'd1381
      10'd46   : in_data <= 14'h0d96; // 'd3478
      10'd47   : in_data <= 14'h1222; // 'd4642
      10'd48   : in_data <= 14'h0ddc; // 'd3548
      10'd49   : in_data <= 14'h0f95; // 'd3989
      10'd50   : in_data <= 14'h00c4; // 'd196
      10'd51   : in_data <= 14'h08d1; // 'd2257
      10'd52   : in_data <= 14'h1319; // 'd4889
      10'd53   : in_data <= 14'h0070; // 'd112
      10'd54   : in_data <= 14'h12bb; // 'd4795
      10'd55   : in_data <= 14'h0866; // 'd2150
      10'd56   : in_data <= 14'h1070; // 'd4208
      10'd57   : in_data <= 14'h0efb; // 'd3835
      10'd58   : in_data <= 14'h12b9; // 'd4793
      10'd59   : in_data <= 14'h1115; // 'd4373
      10'd60   : in_data <= 14'h03dc; // 'd988
      10'd61   : in_data <= 14'h06a6; // 'd1702
      10'd62   : in_data <= 14'h0f52; // 'd3922
      10'd63   : in_data <= 14'h08d5; // 'd2261
      10'd64   : in_data <= 14'h0f0e; // 'd3854
      10'd65   : in_data <= 14'h0474; // 'd1140
      10'd66   : in_data <= 14'h0af2; // 'd2802
      10'd67   : in_data <= 14'h01f2; // 'd498
      10'd68   : in_data <= 14'h0993; // 'd2451
      10'd69   : in_data <= 14'h0056; // 'd86
      10'd70   : in_data <= 14'h0b34; // 'd2868
      10'd71   : in_data <= 14'h1248; // 'd4680
      10'd72   : in_data <= 14'h0149; // 'd329
      10'd73   : in_data <= 14'h0f01; // 'd3841
      10'd74   : in_data <= 14'h0ea2; // 'd3746
      10'd75   : in_data <= 14'h07e4; // 'd2020
      10'd76   : in_data <= 14'h0cee; // 'd3310
      10'd77   : in_data <= 14'h128a; // 'd4746
      10'd78   : in_data <= 14'h0bf7; // 'd3063
      10'd79   : in_data <= 14'h02e7; // 'd743
      10'd80   : in_data <= 14'h03ad; // 'd941
      10'd81   : in_data <= 14'h0952; // 'd2386
      10'd82   : in_data <= 14'h080f; // 'd2063
      10'd83   : in_data <= 14'h0296; // 'd662
      10'd84   : in_data <= 14'h029b; // 'd667
      10'd85   : in_data <= 14'h078c; // 'd1932
      10'd86   : in_data <= 14'h1041; // 'd4161
      10'd87   : in_data <= 14'h0749; // 'd1865
      10'd88   : in_data <= 14'h128f; // 'd4751
      10'd89   : in_data <= 14'h0aa8; // 'd2728
      10'd90   : in_data <= 14'h0c69; // 'd3177
      10'd91   : in_data <= 14'h0389; // 'd905
      10'd92   : in_data <= 14'h05dd; // 'd1501
      10'd93   : in_data <= 14'h06c9; // 'd1737
      10'd94   : in_data <= 14'h00ea; // 'd234
      10'd95   : in_data <= 14'h0985; // 'd2437
      10'd96   : in_data <= 14'h0327; // 'd807
      10'd97   : in_data <= 14'h10c1; // 'd4289
      10'd98   : in_data <= 14'h0d2c; // 'd3372
      10'd99   : in_data <= 14'h1374; // 'd4980
      10'd100  : in_data <= 14'h06ab; // 'd1707
      10'd101  : in_data <= 14'h113a; // 'd4410
      10'd102  : in_data <= 14'h03ea; // 'd1002
      10'd103  : in_data <= 14'h07fc; // 'd2044
      10'd104  : in_data <= 14'h0e03; // 'd3587
      10'd105  : in_data <= 14'h0dd0; // 'd3536
      10'd106  : in_data <= 14'h05b0; // 'd1456
      10'd107  : in_data <= 14'h0048; // 'd72
      10'd108  : in_data <= 14'h12a2; // 'd4770
      10'd109  : in_data <= 14'h1385; // 'd4997
      10'd110  : in_data <= 14'h06df; // 'd1759
      10'd111  : in_data <= 14'h1041; // 'd4161
      10'd112  : in_data <= 14'h0a09; // 'd2569
      10'd113  : in_data <= 14'h1297; // 'd4759
      10'd114  : in_data <= 14'h019d; // 'd413
      10'd115  : in_data <= 14'h069b; // 'd1691
      10'd116  : in_data <= 14'h03d5; // 'd981
      10'd117  : in_data <= 14'h114c; // 'd4428
      10'd118  : in_data <= 14'h112d; // 'd4397
      10'd119  : in_data <= 14'h0d88; // 'd3464
      10'd120  : in_data <= 14'h0f29; // 'd3881
      10'd121  : in_data <= 14'h0740; // 'd1856
      10'd122  : in_data <= 14'h02dd; // 'd733
      10'd123  : in_data <= 14'h004f; // 'd79
      10'd124  : in_data <= 14'h07e3; // 'd2019
      10'd125  : in_data <= 14'h0ea6; // 'd3750
      10'd126  : in_data <= 14'h0ddd; // 'd3549
      10'd127  : in_data <= 14'h11db; // 'd4571
      10'd128  : in_data <= 14'h0474; // 'd1140
      10'd129  : in_data <= 14'h1377; // 'd4983
      10'd130  : in_data <= 14'h050e; // 'd1294
      10'd131  : in_data <= 14'h0df1; // 'd3569
      10'd132  : in_data <= 14'h1150; // 'd4432
      10'd133  : in_data <= 14'h0a9c; // 'd2716
      10'd134  : in_data <= 14'h04b4; // 'd1204
      10'd135  : in_data <= 14'h0a80; // 'd2688
      10'd136  : in_data <= 14'h0e88; // 'd3720
      10'd137  : in_data <= 14'h10ba; // 'd4282
      10'd138  : in_data <= 14'h0f64; // 'd3940
      10'd139  : in_data <= 14'h10d8; // 'd4312
      10'd140  : in_data <= 14'h0e54; // 'd3668
      10'd141  : in_data <= 14'h03e2; // 'd994
      10'd142  : in_data <= 14'h0e08; // 'd3592
      10'd143  : in_data <= 14'h0781; // 'd1921
      10'd144  : in_data <= 14'h1333; // 'd4915
      10'd145  : in_data <= 14'h01ea; // 'd490
      10'd146  : in_data <= 14'h042c; // 'd1068
      10'd147  : in_data <= 14'h05cc; // 'd1484
      10'd148  : in_data <= 14'h1268; // 'd4712
      10'd149  : in_data <= 14'h0dfe; // 'd3582
      10'd150  : in_data <= 14'h0e28; // 'd3624
      10'd151  : in_data <= 14'h00a4; // 'd164
      10'd152  : in_data <= 14'h008c; // 'd140
      10'd153  : in_data <= 14'h081a; // 'd2074
      10'd154  : in_data <= 14'h058b; // 'd1419
      10'd155  : in_data <= 14'h116e; // 'd4462
      10'd156  : in_data <= 14'h116b; // 'd4459
      10'd157  : in_data <= 14'h0a87; // 'd2695
      10'd158  : in_data <= 14'h0a26; // 'd2598
      10'd159  : in_data <= 14'h0703; // 'd1795
      10'd160  : in_data <= 14'h1330; // 'd4912
      10'd161  : in_data <= 14'h00f3; // 'd243
      10'd162  : in_data <= 14'h1234; // 'd4660
      10'd163  : in_data <= 14'h05b0; // 'd1456
      10'd164  : in_data <= 14'h04fa; // 'd1274
      10'd165  : in_data <= 14'h0853; // 'd2131
      10'd166  : in_data <= 14'h0af7; // 'd2807
      10'd167  : in_data <= 14'h11e9; // 'd4585
      10'd168  : in_data <= 14'h1424; // 'd5156
      10'd169  : in_data <= 14'h0c11; // 'd3089
      10'd170  : in_data <= 14'h13c6; // 'd5062
      10'd171  : in_data <= 14'h0bf7; // 'd3063
      10'd172  : in_data <= 14'h05ac; // 'd1452
      10'd173  : in_data <= 14'h028d; // 'd653
      10'd174  : in_data <= 14'h0f0e; // 'd3854
      10'd175  : in_data <= 14'h10b1; // 'd4273
      10'd176  : in_data <= 14'h004f; // 'd79
      10'd177  : in_data <= 14'h0775; // 'd1909
      10'd178  : in_data <= 14'h0940; // 'd2368
      10'd179  : in_data <= 14'h0635; // 'd1589
      10'd180  : in_data <= 14'h11fd; // 'd4605
      10'd181  : in_data <= 14'h0453; // 'd1107
      10'd182  : in_data <= 14'h07c2; // 'd1986
      10'd183  : in_data <= 14'h0f9c; // 'd3996
      10'd184  : in_data <= 14'h06ff; // 'd1791
      10'd185  : in_data <= 14'h0867; // 'd2151
      10'd186  : in_data <= 14'h0050; // 'd80
      10'd187  : in_data <= 14'h1356; // 'd4950
      10'd188  : in_data <= 14'h0c11; // 'd3089
      10'd189  : in_data <= 14'h1414; // 'd5140
      10'd190  : in_data <= 14'h0442; // 'd1090
      10'd191  : in_data <= 14'h041e; // 'd1054
      10'd192  : in_data <= 14'h06b8; // 'd1720
      10'd193  : in_data <= 14'h0d78; // 'd3448
      10'd194  : in_data <= 14'h0819; // 'd2073
      10'd195  : in_data <= 14'h0176; // 'd374
      10'd196  : in_data <= 14'h0e80; // 'd3712
      10'd197  : in_data <= 14'h04fd; // 'd1277
      10'd198  : in_data <= 14'h0085; // 'd133
      10'd199  : in_data <= 14'h0bf2; // 'd3058
      10'd200  : in_data <= 14'h09b4; // 'd2484
      10'd201  : in_data <= 14'h136c; // 'd4972
      10'd202  : in_data <= 14'h05a1; // 'd1441
      10'd203  : in_data <= 14'h04bb; // 'd1211
      10'd204  : in_data <= 14'h0e59; // 'd3673
      10'd205  : in_data <= 14'h09ea; // 'd2538
      10'd206  : in_data <= 14'h1255; // 'd4693
      10'd207  : in_data <= 14'h068e; // 'd1678
      10'd208  : in_data <= 14'h043c; // 'd1084
      10'd209  : in_data <= 14'h10a4; // 'd4260
      10'd210  : in_data <= 14'h007e; // 'd126
      10'd211  : in_data <= 14'h0422; // 'd1058
      10'd212  : in_data <= 14'h140f; // 'd5135
      10'd213  : in_data <= 14'h066a; // 'd1642
      10'd214  : in_data <= 14'h0097; // 'd151
      10'd215  : in_data <= 14'h00bc; // 'd188
      10'd216  : in_data <= 14'h0c92; // 'd3218
      10'd217  : in_data <= 14'h0bc0; // 'd3008
      10'd218  : in_data <= 14'h10c2; // 'd4290
      10'd219  : in_data <= 14'h0e1b; // 'd3611
      10'd220  : in_data <= 14'h03ac; // 'd940
      10'd221  : in_data <= 14'h0877; // 'd2167
      10'd222  : in_data <= 14'h11bc; // 'd4540
      10'd223  : in_data <= 14'h04c4; // 'd1220
      10'd224  : in_data <= 14'h02b8; // 'd696
      10'd225  : in_data <= 14'h141e; // 'd5150
      10'd226  : in_data <= 14'h13e1; // 'd5089
      10'd227  : in_data <= 14'h0e56; // 'd3670
      10'd228  : in_data <= 14'h12fb; // 'd4859
      10'd229  : in_data <= 14'h05eb; // 'd1515
      10'd230  : in_data <= 14'h0d77; // 'd3447
      10'd231  : in_data <= 14'h0322; // 'd802
      10'd232  : in_data <= 14'h059a; // 'd1434
      10'd233  : in_data <= 14'h03ca; // 'd970
      10'd234  : in_data <= 14'h116d; // 'd4461
      10'd235  : in_data <= 14'h0498; // 'd1176
      10'd236  : in_data <= 14'h021f; // 'd543
      10'd237  : in_data <= 14'h0067; // 'd103
      10'd238  : in_data <= 14'h03a1; // 'd929
      10'd239  : in_data <= 14'h10b0; // 'd4272
      10'd240  : in_data <= 14'h0f5e; // 'd3934
      10'd241  : in_data <= 14'h1039; // 'd4153
      10'd242  : in_data <= 14'h0054; // 'd84
      10'd243  : in_data <= 14'h01a9; // 'd425
      10'd244  : in_data <= 14'h045a; // 'd1114
      10'd245  : in_data <= 14'h08ef; // 'd2287
      10'd246  : in_data <= 14'h091a; // 'd2330
      10'd247  : in_data <= 14'h062a; // 'd1578
      10'd248  : in_data <= 14'h01cd; // 'd461
      10'd249  : in_data <= 14'h0938; // 'd2360
      10'd250  : in_data <= 14'h0041; // 'd65
      10'd251  : in_data <= 14'h112b; // 'd4395
      10'd252  : in_data <= 14'h0710; // 'd1808
      10'd253  : in_data <= 14'h05af; // 'd1455
      10'd254  : in_data <= 14'h077b; // 'd1915
      10'd255  : in_data <= 14'h0404; // 'd1028
      10'd256  : in_data <= 14'h06fc; // 'd1788
      10'd257  : in_data <= 14'h0db8; // 'd3512
      10'd258  : in_data <= 14'h03c5; // 'd965
      10'd259  : in_data <= 14'h082e; // 'd2094
      10'd260  : in_data <= 14'h02bb; // 'd699
      10'd261  : in_data <= 14'h043c; // 'd1084
      10'd262  : in_data <= 14'h0ea8; // 'd3752
      10'd263  : in_data <= 14'h04f8; // 'd1272
      10'd264  : in_data <= 14'h0c5b; // 'd3163
      10'd265  : in_data <= 14'h020c; // 'd524
      10'd266  : in_data <= 14'h024a; // 'd586
      10'd267  : in_data <= 14'h1087; // 'd4231
      10'd268  : in_data <= 14'h0e67; // 'd3687
      10'd269  : in_data <= 14'h0e55; // 'd3669
      10'd270  : in_data <= 14'h023e; // 'd574
      10'd271  : in_data <= 14'h1039; // 'd4153
      10'd272  : in_data <= 14'h0e5c; // 'd3676
      10'd273  : in_data <= 14'h0056; // 'd86
      10'd274  : in_data <= 14'h0187; // 'd391
      10'd275  : in_data <= 14'h005d; // 'd93
      10'd276  : in_data <= 14'h1193; // 'd4499
      10'd277  : in_data <= 14'h0ddf; // 'd3551
      10'd278  : in_data <= 14'h11b4; // 'd4532
      10'd279  : in_data <= 14'h0812; // 'd2066
      10'd280  : in_data <= 14'h0c08; // 'd3080
      10'd281  : in_data <= 14'h129a; // 'd4762
      10'd282  : in_data <= 14'h0956; // 'd2390
      10'd283  : in_data <= 14'h06a0; // 'd1696
      10'd284  : in_data <= 14'h03fd; // 'd1021
      10'd285  : in_data <= 14'h0cc8; // 'd3272
      10'd286  : in_data <= 14'h0c16; // 'd3094
      10'd287  : in_data <= 14'h09a8; // 'd2472
      10'd288  : in_data <= 14'h0fa5; // 'd4005
      10'd289  : in_data <= 14'h13b3; // 'd5043
      10'd290  : in_data <= 14'h0c43; // 'd3139
      10'd291  : in_data <= 14'h1378; // 'd4984
      10'd292  : in_data <= 14'h0103; // 'd259
      10'd293  : in_data <= 14'h13dc; // 'd5084
      10'd294  : in_data <= 14'h1128; // 'd4392
      10'd295  : in_data <= 14'h0508; // 'd1288
      10'd296  : in_data <= 14'h13fd; // 'd5117
      10'd297  : in_data <= 14'h1096; // 'd4246
      10'd298  : in_data <= 14'h1180; // 'd4480
      10'd299  : in_data <= 14'h0714; // 'd1812
      10'd300  : in_data <= 14'h0dfa; // 'd3578
      10'd301  : in_data <= 14'h0c89; // 'd3209
      10'd302  : in_data <= 14'h0f2c; // 'd3884
      10'd303  : in_data <= 14'h009c; // 'd156
      10'd304  : in_data <= 14'h10ec; // 'd4332
      10'd305  : in_data <= 14'h0a13; // 'd2579
      10'd306  : in_data <= 14'h098a; // 'd2442
      10'd307  : in_data <= 14'h04ff; // 'd1279
      10'd308  : in_data <= 14'h1175; // 'd4469
      10'd309  : in_data <= 14'h115f; // 'd4447
      10'd310  : in_data <= 14'h0069; // 'd105
      10'd311  : in_data <= 14'h131f; // 'd4895
      10'd312  : in_data <= 14'h138b; // 'd5003
      10'd313  : in_data <= 14'h0ba0; // 'd2976
      10'd314  : in_data <= 14'h0a37; // 'd2615
      10'd315  : in_data <= 14'h0e34; // 'd3636
      10'd316  : in_data <= 14'h1360; // 'd4960
      10'd317  : in_data <= 14'h1087; // 'd4231
      10'd318  : in_data <= 14'h0f38; // 'd3896
      10'd319  : in_data <= 14'h0f7f; // 'd3967
      10'd320  : in_data <= 14'h071f; // 'd1823
      10'd321  : in_data <= 14'h0750; // 'd1872
      10'd322  : in_data <= 14'h00bf; // 'd191
      10'd323  : in_data <= 14'h02b5; // 'd693
      10'd324  : in_data <= 14'h0247; // 'd583
      10'd325  : in_data <= 14'h0138; // 'd312
      10'd326  : in_data <= 14'h097a; // 'd2426
      10'd327  : in_data <= 14'h0c89; // 'd3209
      10'd328  : in_data <= 14'h0149; // 'd329
      10'd329  : in_data <= 14'h0e12; // 'd3602
      10'd330  : in_data <= 14'h1058; // 'd4184
      10'd331  : in_data <= 14'h0df2; // 'd3570
      10'd332  : in_data <= 14'h00ea; // 'd234
      10'd333  : in_data <= 14'h03f7; // 'd1015
      10'd334  : in_data <= 14'h1126; // 'd4390
      10'd335  : in_data <= 14'h0c63; // 'd3171
      10'd336  : in_data <= 14'h115d; // 'd4445
      10'd337  : in_data <= 14'h0dcc; // 'd3532
      10'd338  : in_data <= 14'h07d9; // 'd2009
      10'd339  : in_data <= 14'h0e13; // 'd3603
      10'd340  : in_data <= 14'h04b4; // 'd1204
      10'd341  : in_data <= 14'h0e6c; // 'd3692
      10'd342  : in_data <= 14'h10ea; // 'd4330
      10'd343  : in_data <= 14'h1103; // 'd4355
      10'd344  : in_data <= 14'h0195; // 'd405
      10'd345  : in_data <= 14'h0612; // 'd1554
      10'd346  : in_data <= 14'h09cb; // 'd2507
      10'd347  : in_data <= 14'h1221; // 'd4641
      10'd348  : in_data <= 14'h0609; // 'd1545
      10'd349  : in_data <= 14'h0eb8; // 'd3768
      10'd350  : in_data <= 14'h0f78; // 'd3960
      10'd351  : in_data <= 14'h02ac; // 'd684
      10'd352  : in_data <= 14'h0ac7; // 'd2759
      10'd353  : in_data <= 14'h0224; // 'd548
      10'd354  : in_data <= 14'h003a; // 'd58
      10'd355  : in_data <= 14'h0b12; // 'd2834
      10'd356  : in_data <= 14'h0582; // 'd1410
      10'd357  : in_data <= 14'h0ad3; // 'd2771
      10'd358  : in_data <= 14'h008f; // 'd143
      10'd359  : in_data <= 14'h0fbd; // 'd4029
      10'd360  : in_data <= 14'h0c4e; // 'd3150
      10'd361  : in_data <= 14'h0a74; // 'd2676
      10'd362  : in_data <= 14'h0671; // 'd1649
      10'd363  : in_data <= 14'h0daf; // 'd3503
      10'd364  : in_data <= 14'h037c; // 'd892
      10'd365  : in_data <= 14'h018b; // 'd395
      10'd366  : in_data <= 14'h0566; // 'd1382
      10'd367  : in_data <= 14'h12e0; // 'd4832
      10'd368  : in_data <= 14'h0f6c; // 'd3948
      10'd369  : in_data <= 14'h0f8b; // 'd3979
      10'd370  : in_data <= 14'h13f1; // 'd5105
      10'd371  : in_data <= 14'h103b; // 'd4155
      10'd372  : in_data <= 14'h08e8; // 'd2280
      10'd373  : in_data <= 14'h124b; // 'd4683
      10'd374  : in_data <= 14'h0ce7; // 'd3303
      10'd375  : in_data <= 14'h0408; // 'd1032
      10'd376  : in_data <= 14'h11c4; // 'd4548
      10'd377  : in_data <= 14'h0e31; // 'd3633
      10'd378  : in_data <= 14'h0b1f; // 'd2847
      10'd379  : in_data <= 14'h0906; // 'd2310
      10'd380  : in_data <= 14'h066e; // 'd1646
      10'd381  : in_data <= 14'h055b; // 'd1371
      10'd382  : in_data <= 14'h0b7c; // 'd2940
      10'd383  : in_data <= 14'h0d79; // 'd3449
      10'd384  : in_data <= 14'h0ae5; // 'd2789
      10'd385  : in_data <= 14'h099f; // 'd2463
      10'd386  : in_data <= 14'h06fc; // 'd1788
      10'd387  : in_data <= 14'h0ab2; // 'd2738
      10'd388  : in_data <= 14'h099c; // 'd2460
      10'd389  : in_data <= 14'h1186; // 'd4486
      10'd390  : in_data <= 14'h02bb; // 'd699
      10'd391  : in_data <= 14'h07cf; // 'd1999
      10'd392  : in_data <= 14'h047e; // 'd1150
      10'd393  : in_data <= 14'h0349; // 'd841
      10'd394  : in_data <= 14'h0a30; // 'd2608
      10'd395  : in_data <= 14'h1424; // 'd5156
      10'd396  : in_data <= 14'h0e21; // 'd3617
      10'd397  : in_data <= 14'h0ea0; // 'd3744
      10'd398  : in_data <= 14'h06cd; // 'd1741
      10'd399  : in_data <= 14'h061d; // 'd1565
      10'd400  : in_data <= 14'h0b84; // 'd2948
      10'd401  : in_data <= 14'h04ef; // 'd1263
      10'd402  : in_data <= 14'h078f; // 'd1935
      10'd403  : in_data <= 14'h11fc; // 'd4604
      10'd404  : in_data <= 14'h0121; // 'd289
      10'd405  : in_data <= 14'h113f; // 'd4415
      10'd406  : in_data <= 14'h111d; // 'd4381
      10'd407  : in_data <= 14'h03b2; // 'd946
      10'd408  : in_data <= 14'h1268; // 'd4712
      10'd409  : in_data <= 14'h0005; // 'd5
      10'd410  : in_data <= 14'h00e3; // 'd227
      10'd411  : in_data <= 14'h1007; // 'd4103
      10'd412  : in_data <= 14'h0c37; // 'd3127
      10'd413  : in_data <= 14'h01bf; // 'd447
      10'd414  : in_data <= 14'h00bf; // 'd191
      10'd415  : in_data <= 14'h0963; // 'd2403
      10'd416  : in_data <= 14'h110b; // 'd4363
      10'd417  : in_data <= 14'h0f89; // 'd3977
      10'd418  : in_data <= 14'h0ce3; // 'd3299
      10'd419  : in_data <= 14'h002c; // 'd44
      10'd420  : in_data <= 14'h13cd; // 'd5069
      10'd421  : in_data <= 14'h0f43; // 'd3907
      10'd422  : in_data <= 14'h049a; // 'd1178
      10'd423  : in_data <= 14'h0b93; // 'd2963
      10'd424  : in_data <= 14'h1211; // 'd4625
      10'd425  : in_data <= 14'h076f; // 'd1903
      10'd426  : in_data <= 14'h017f; // 'd383
      10'd427  : in_data <= 14'h0506; // 'd1286
      10'd428  : in_data <= 14'h0164; // 'd356
      10'd429  : in_data <= 14'h0e31; // 'd3633
      10'd430  : in_data <= 14'h0e79; // 'd3705
      10'd431  : in_data <= 14'h13e9; // 'd5097
      10'd432  : in_data <= 14'h0636; // 'd1590
      10'd433  : in_data <= 14'h1246; // 'd4678
      10'd434  : in_data <= 14'h0cc2; // 'd3266
      10'd435  : in_data <= 14'h010c; // 'd268
      10'd436  : in_data <= 14'h140e; // 'd5134
      10'd437  : in_data <= 14'h032f; // 'd815
      10'd438  : in_data <= 14'h1390; // 'd5008
      10'd439  : in_data <= 14'h067f; // 'd1663
      10'd440  : in_data <= 14'h0369; // 'd873
      10'd441  : in_data <= 14'h0bb5; // 'd2997
      10'd442  : in_data <= 14'h0fa6; // 'd4006
      10'd443  : in_data <= 14'h1184; // 'd4484
      10'd444  : in_data <= 14'h00f7; // 'd247
      10'd445  : in_data <= 14'h0196; // 'd406
      10'd446  : in_data <= 14'h046b; // 'd1131
      10'd447  : in_data <= 14'h0159; // 'd345
      10'd448  : in_data <= 14'h10e4; // 'd4324
      10'd449  : in_data <= 14'h12c7; // 'd4807
      10'd450  : in_data <= 14'h06d7; // 'd1751
      10'd451  : in_data <= 14'h11d6; // 'd4566
      10'd452  : in_data <= 14'h0a44; // 'd2628
      10'd453  : in_data <= 14'h047e; // 'd1150
      10'd454  : in_data <= 14'h0d6d; // 'd3437
      10'd455  : in_data <= 14'h052e; // 'd1326
      10'd456  : in_data <= 14'h08ab; // 'd2219
      10'd457  : in_data <= 14'h13ce; // 'd5070
      10'd458  : in_data <= 14'h03ee; // 'd1006
      10'd459  : in_data <= 14'h025a; // 'd602
      10'd460  : in_data <= 14'h138a; // 'd5002
      10'd461  : in_data <= 14'h07df; // 'd2015
      10'd462  : in_data <= 14'h0908; // 'd2312
      10'd463  : in_data <= 14'h0b10; // 'd2832
      10'd464  : in_data <= 14'h11cd; // 'd4557
      10'd465  : in_data <= 14'h0cbe; // 'd3262
      10'd466  : in_data <= 14'h1000; // 'd4096
      10'd467  : in_data <= 14'h0cb2; // 'd3250
      10'd468  : in_data <= 14'h0106; // 'd262
      10'd469  : in_data <= 14'h0db4; // 'd3508
      10'd470  : in_data <= 14'h0f7a; // 'd3962
      10'd471  : in_data <= 14'h0f1b; // 'd3867
      10'd472  : in_data <= 14'h0a3d; // 'd2621
      10'd473  : in_data <= 14'h0639; // 'd1593
      10'd474  : in_data <= 14'h063f; // 'd1599
      10'd475  : in_data <= 14'h0a71; // 'd2673
      10'd476  : in_data <= 14'h0d2a; // 'd3370
      10'd477  : in_data <= 14'h0b89; // 'd2953
      10'd478  : in_data <= 14'h06e6; // 'd1766
      10'd479  : in_data <= 14'h0325; // 'd805
      10'd480  : in_data <= 14'h1373; // 'd4979
      10'd481  : in_data <= 14'h0eb6; // 'd3766
      10'd482  : in_data <= 14'h09a6; // 'd2470
      10'd483  : in_data <= 14'h0177; // 'd375
      10'd484  : in_data <= 14'h0ee1; // 'd3809
      10'd485  : in_data <= 14'h09ab; // 'd2475
      10'd486  : in_data <= 14'h0288; // 'd648
      10'd487  : in_data <= 14'h1055; // 'd4181
      10'd488  : in_data <= 14'h07bf; // 'd1983
      10'd489  : in_data <= 14'h0bf5; // 'd3061
      10'd490  : in_data <= 14'h0255; // 'd597
      10'd491  : in_data <= 14'h01f0; // 'd496
      10'd492  : in_data <= 14'h0553; // 'd1363
      10'd493  : in_data <= 14'h0d7b; // 'd3451
      10'd494  : in_data <= 14'h050f; // 'd1295
      10'd495  : in_data <= 14'h0d07; // 'd3335
      10'd496  : in_data <= 14'h0e0a; // 'd3594
      10'd497  : in_data <= 14'h1147; // 'd4423
      10'd498  : in_data <= 14'h0dc9; // 'd3529
      10'd499  : in_data <= 14'h0d67; // 'd3431
      10'd500  : in_data <= 14'h0cd3; // 'd3283
      10'd501  : in_data <= 14'h07bb; // 'd1979
      10'd502  : in_data <= 14'h106e; // 'd4206
      10'd503  : in_data <= 14'h0273; // 'd627
      10'd504  : in_data <= 14'h0a7c; // 'd2684
      10'd505  : in_data <= 14'h031a; // 'd794
      10'd506  : in_data <= 14'h12a4; // 'd4772
      10'd507  : in_data <= 14'h0c9f; // 'd3231
      10'd508  : in_data <= 14'h0344; // 'd836
      10'd509  : in_data <= 14'h0826; // 'd2086
      10'd510  : in_data <= 14'h0b78; // 'd2936
      10'd511  : in_data <= 14'h0fae; // 'd4014
      10'd512  : in_data <= 14'h00f6; // 'd246
      10'd513  : in_data <= 14'h11d9; // 'd4569
      10'd514  : in_data <= 14'h13e0; // 'd5088
      10'd515  : in_data <= 14'h1037; // 'd4151
      10'd516  : in_data <= 14'h1315; // 'd4885
      10'd517  : in_data <= 14'h052c; // 'd1324
      10'd518  : in_data <= 14'h0e1c; // 'd3612
      10'd519  : in_data <= 14'h12cf; // 'd4815
      10'd520  : in_data <= 14'h1022; // 'd4130
      10'd521  : in_data <= 14'h10ad; // 'd4269
      10'd522  : in_data <= 14'h0d99; // 'd3481
      10'd523  : in_data <= 14'h101b; // 'd4123
      10'd524  : in_data <= 14'h104d; // 'd4173
      10'd525  : in_data <= 14'h0843; // 'd2115
      10'd526  : in_data <= 14'h0a7e; // 'd2686
      10'd527  : in_data <= 14'h0d72; // 'd3442
      10'd528  : in_data <= 14'h0891; // 'd2193
      10'd529  : in_data <= 14'h05a8; // 'd1448
      10'd530  : in_data <= 14'h12d4; // 'd4820
      10'd531  : in_data <= 14'h0305; // 'd773
      10'd532  : in_data <= 14'h06bd; // 'd1725
      10'd533  : in_data <= 14'h0fba; // 'd4026
      10'd534  : in_data <= 14'h0538; // 'd1336
      10'd535  : in_data <= 14'h0a0e; // 'd2574
      10'd536  : in_data <= 14'h0d3e; // 'd3390
      10'd537  : in_data <= 14'h07ed; // 'd2029
      10'd538  : in_data <= 14'h0f90; // 'd3984
      10'd539  : in_data <= 14'h141e; // 'd5150
      10'd540  : in_data <= 14'h107e; // 'd4222
      10'd541  : in_data <= 14'h08c7; // 'd2247
      10'd542  : in_data <= 14'h02ae; // 'd686
      10'd543  : in_data <= 14'h1084; // 'd4228
      10'd544  : in_data <= 14'h0ea1; // 'd3745
      10'd545  : in_data <= 14'h0c41; // 'd3137
      10'd546  : in_data <= 14'h1408; // 'd5128
      10'd547  : in_data <= 14'h0143; // 'd323
      10'd548  : in_data <= 14'h0b99; // 'd2969
      10'd549  : in_data <= 14'h0889; // 'd2185
      10'd550  : in_data <= 14'h05d3; // 'd1491
      10'd551  : in_data <= 14'h08c3; // 'd2243
      10'd552  : in_data <= 14'h03d5; // 'd981
      10'd553  : in_data <= 14'h01bb; // 'd443
      10'd554  : in_data <= 14'h1330; // 'd4912
      10'd555  : in_data <= 14'h0a2d; // 'd2605
      10'd556  : in_data <= 14'h0df6; // 'd3574
      10'd557  : in_data <= 14'h06fd; // 'd1789
      10'd558  : in_data <= 14'h0677; // 'd1655
      10'd559  : in_data <= 14'h0e57; // 'd3671
      10'd560  : in_data <= 14'h0ed2; // 'd3794
      10'd561  : in_data <= 14'h0285; // 'd645
      10'd562  : in_data <= 14'h064b; // 'd1611
      10'd563  : in_data <= 14'h0f46; // 'd3910
      10'd564  : in_data <= 14'h037b; // 'd891
      10'd565  : in_data <= 14'h02d6; // 'd726
      10'd566  : in_data <= 14'h0521; // 'd1313
      10'd567  : in_data <= 14'h0b40; // 'd2880
      10'd568  : in_data <= 14'h139e; // 'd5022
      10'd569  : in_data <= 14'h12e5; // 'd4837
      10'd570  : in_data <= 14'h0d6d; // 'd3437
      10'd571  : in_data <= 14'h0b38; // 'd2872
      10'd572  : in_data <= 14'h087b; // 'd2171
      10'd573  : in_data <= 14'h0414; // 'd1044
      10'd574  : in_data <= 14'h0dd3; // 'd3539
      10'd575  : in_data <= 14'h1204; // 'd4612
      10'd576  : in_data <= 14'h0ff4; // 'd4084
      10'd577  : in_data <= 14'h0a3e; // 'd2622
      10'd578  : in_data <= 14'h08a7; // 'd2215
      10'd579  : in_data <= 14'h008a; // 'd138
      10'd580  : in_data <= 14'h02b8; // 'd696
      10'd581  : in_data <= 14'h099f; // 'd2463
      10'd582  : in_data <= 14'h0ef6; // 'd3830
      10'd583  : in_data <= 14'h00e1; // 'd225
      10'd584  : in_data <= 14'h0890; // 'd2192
      10'd585  : in_data <= 14'h0e42; // 'd3650
      10'd586  : in_data <= 14'h100f; // 'd4111
      10'd587  : in_data <= 14'h090e; // 'd2318
      10'd588  : in_data <= 14'h03b1; // 'd945
      10'd589  : in_data <= 14'h0364; // 'd868
      10'd590  : in_data <= 14'h0bbe; // 'd3006
      10'd591  : in_data <= 14'h12a4; // 'd4772
      10'd592  : in_data <= 14'h0936; // 'd2358
      10'd593  : in_data <= 14'h0067; // 'd103
      10'd594  : in_data <= 14'h0600; // 'd1536
      10'd595  : in_data <= 14'h080b; // 'd2059
      10'd596  : in_data <= 14'h01dc; // 'd476
      10'd597  : in_data <= 14'h0a3d; // 'd2621
      10'd598  : in_data <= 14'h12da; // 'd4826
      10'd599  : in_data <= 14'h13fb; // 'd5115
      10'd600  : in_data <= 14'h002a; // 'd42
      10'd601  : in_data <= 14'h0d77; // 'd3447
      10'd602  : in_data <= 14'h072a; // 'd1834
      10'd603  : in_data <= 14'h0e49; // 'd3657
      10'd604  : in_data <= 14'h0e5a; // 'd3674
      10'd605  : in_data <= 14'h0f19; // 'd3865
      10'd606  : in_data <= 14'h040f; // 'd1039
      10'd607  : in_data <= 14'h07e6; // 'd2022
      10'd608  : in_data <= 14'h0c50; // 'd3152
      10'd609  : in_data <= 14'h0480; // 'd1152
      10'd610  : in_data <= 14'h12ec; // 'd4844
      10'd611  : in_data <= 14'h0cc5; // 'd3269
      10'd612  : in_data <= 14'h0a36; // 'd2614
      10'd613  : in_data <= 14'h1173; // 'd4467
      10'd614  : in_data <= 14'h0192; // 'd402
      10'd615  : in_data <= 14'h042a; // 'd1066
      10'd616  : in_data <= 14'h0e11; // 'd3601
      10'd617  : in_data <= 14'h0cc6; // 'd3270
      10'd618  : in_data <= 14'h0f18; // 'd3864
      10'd619  : in_data <= 14'h0b7a; // 'd2938
      10'd620  : in_data <= 14'h0152; // 'd338
      10'd621  : in_data <= 14'h0af1; // 'd2801
      10'd622  : in_data <= 14'h0e98; // 'd3736
      10'd623  : in_data <= 14'h0618; // 'd1560
      10'd624  : in_data <= 14'h0196; // 'd406
      10'd625  : in_data <= 14'h0182; // 'd386
      10'd626  : in_data <= 14'h1298; // 'd4760
      10'd627  : in_data <= 14'h126e; // 'd4718
      10'd628  : in_data <= 14'h05d4; // 'd1492
      10'd629  : in_data <= 14'h0ba7; // 'd2983
      10'd630  : in_data <= 14'h0fa8; // 'd4008
      10'd631  : in_data <= 14'h0049; // 'd73
      10'd632  : in_data <= 14'h0562; // 'd1378
      10'd633  : in_data <= 14'h125d; // 'd4701
      10'd634  : in_data <= 14'h0f68; // 'd3944
      10'd635  : in_data <= 14'h0f54; // 'd3924
      10'd636  : in_data <= 14'h1402; // 'd5122
      10'd637  : in_data <= 14'h0526; // 'd1318
      10'd638  : in_data <= 14'h0495; // 'd1173
      10'd639  : in_data <= 14'h0731; // 'd1841
      10'd640  : in_data <= 14'h0d2f; // 'd3375
      10'd641  : in_data <= 14'h131a; // 'd4890
      10'd642  : in_data <= 14'h0825; // 'd2085
      10'd643  : in_data <= 14'h024d; // 'd589
      10'd644  : in_data <= 14'h1066; // 'd4198
      10'd645  : in_data <= 14'h0ad1; // 'd2769
      10'd646  : in_data <= 14'h05ad; // 'd1453
      10'd647  : in_data <= 14'h10eb; // 'd4331
      10'd648  : in_data <= 14'h1398; // 'd5016
      10'd649  : in_data <= 14'h0514; // 'd1300
      10'd650  : in_data <= 14'h0d02; // 'd3330
      10'd651  : in_data <= 14'h0e0b; // 'd3595
      10'd652  : in_data <= 14'h05ce; // 'd1486
      10'd653  : in_data <= 14'h0294; // 'd660
      10'd654  : in_data <= 14'h0b7d; // 'd2941
      10'd655  : in_data <= 14'h0522; // 'd1314
      10'd656  : in_data <= 14'h0a77; // 'd2679
      10'd657  : in_data <= 14'h0e1a; // 'd3610
      10'd658  : in_data <= 14'h0b12; // 'd2834
      10'd659  : in_data <= 14'h095b; // 'd2395
      10'd660  : in_data <= 14'h023e; // 'd574
      10'd661  : in_data <= 14'h05da; // 'd1498
      10'd662  : in_data <= 14'h0b71; // 'd2929
      10'd663  : in_data <= 14'h07e7; // 'd2023
      10'd664  : in_data <= 14'h0d20; // 'd3360
      10'd665  : in_data <= 14'h0203; // 'd515
      10'd666  : in_data <= 14'h0f0d; // 'd3853
      10'd667  : in_data <= 14'h0c19; // 'd3097
      10'd668  : in_data <= 14'h0fe8; // 'd4072
      10'd669  : in_data <= 14'h0845; // 'd2117
      10'd670  : in_data <= 14'h05d7; // 'd1495
      10'd671  : in_data <= 14'h0234; // 'd564
      10'd672  : in_data <= 14'h053d; // 'd1341
      10'd673  : in_data <= 14'h1184; // 'd4484
      10'd674  : in_data <= 14'h0e42; // 'd3650
      10'd675  : in_data <= 14'h0af7; // 'd2807
      10'd676  : in_data <= 14'h0c20; // 'd3104
      10'd677  : in_data <= 14'h13cc; // 'd5068
      10'd678  : in_data <= 14'h0a5a; // 'd2650
      10'd679  : in_data <= 14'h1424; // 'd5156
      10'd680  : in_data <= 14'h11d2; // 'd4562
      10'd681  : in_data <= 14'h0121; // 'd289
      10'd682  : in_data <= 14'h0a2e; // 'd2606
      10'd683  : in_data <= 14'h064d; // 'd1613
      10'd684  : in_data <= 14'h03ba; // 'd954
      10'd685  : in_data <= 14'h095e; // 'd2398
      10'd686  : in_data <= 14'h10c9; // 'd4297
      10'd687  : in_data <= 14'h1083; // 'd4227
      10'd688  : in_data <= 14'h0ba1; // 'd2977
      10'd689  : in_data <= 14'h0052; // 'd82
      10'd690  : in_data <= 14'h022e; // 'd558
      10'd691  : in_data <= 14'h0eb3; // 'd3763
      10'd692  : in_data <= 14'h13e7; // 'd5095
      10'd693  : in_data <= 14'h0f75; // 'd3957
      10'd694  : in_data <= 14'h06fe; // 'd1790
      10'd695  : in_data <= 14'h03f9; // 'd1017
      10'd696  : in_data <= 14'h05f7; // 'd1527
      10'd697  : in_data <= 14'h0970; // 'd2416
      10'd698  : in_data <= 14'h0d8e; // 'd3470
      10'd699  : in_data <= 14'h006a; // 'd106
      10'd700  : in_data <= 14'h0cb9; // 'd3257
      10'd701  : in_data <= 14'h084a; // 'd2122
      10'd702  : in_data <= 14'h00c2; // 'd194
      10'd703  : in_data <= 14'h108e; // 'd4238
      10'd704  : in_data <= 14'h0874; // 'd2164
      10'd705  : in_data <= 14'h11d0; // 'd4560
      10'd706  : in_data <= 14'h1277; // 'd4727
      10'd707  : in_data <= 14'h0e92; // 'd3730
      10'd708  : in_data <= 14'h0e87; // 'd3719
      10'd709  : in_data <= 14'h0cf7; // 'd3319
      10'd710  : in_data <= 14'h04d1; // 'd1233
      10'd711  : in_data <= 14'h049e; // 'd1182
      10'd712  : in_data <= 14'h0fb9; // 'd4025
      10'd713  : in_data <= 14'h0a7c; // 'd2684
      10'd714  : in_data <= 14'h08ef; // 'd2287
      10'd715  : in_data <= 14'h1180; // 'd4480
      10'd716  : in_data <= 14'h0e20; // 'd3616
      10'd717  : in_data <= 14'h064d; // 'd1613
      10'd718  : in_data <= 14'h0fb8; // 'd4024
      10'd719  : in_data <= 14'h0160; // 'd352
      10'd720  : in_data <= 14'h0f26; // 'd3878
      10'd721  : in_data <= 14'h11f1; // 'd4593
      10'd722  : in_data <= 14'h03e2; // 'd994
      10'd723  : in_data <= 14'h026f; // 'd623
      10'd724  : in_data <= 14'h01a6; // 'd422
      10'd725  : in_data <= 14'h0fcb; // 'd4043
      10'd726  : in_data <= 14'h0b77; // 'd2935
      10'd727  : in_data <= 14'h0761; // 'd1889
      10'd728  : in_data <= 14'h05d6; // 'd1494
      10'd729  : in_data <= 14'h0732; // 'd1842
      10'd730  : in_data <= 14'h0907; // 'd2311
      10'd731  : in_data <= 14'h0288; // 'd648
      10'd732  : in_data <= 14'h13e2; // 'd5090
      10'd733  : in_data <= 14'h0f80; // 'd3968
      10'd734  : in_data <= 14'h131a; // 'd4890
      10'd735  : in_data <= 14'h1234; // 'd4660
      10'd736  : in_data <= 14'h0018; // 'd24
      10'd737  : in_data <= 14'h056a; // 'd1386
      10'd738  : in_data <= 14'h03f7; // 'd1015
      10'd739  : in_data <= 14'h0dda; // 'd3546
      10'd740  : in_data <= 14'h0031; // 'd49
      10'd741  : in_data <= 14'h03a8; // 'd936
      10'd742  : in_data <= 14'h0737; // 'd1847
      10'd743  : in_data <= 14'h106b; // 'd4203
      10'd744  : in_data <= 14'h0c1c; // 'd3100
      10'd745  : in_data <= 14'h0cf1; // 'd3313
      10'd746  : in_data <= 14'h0d15; // 'd3349
      10'd747  : in_data <= 14'h0b0f; // 'd2831
      10'd748  : in_data <= 14'h0546; // 'd1350
      10'd749  : in_data <= 14'h0529; // 'd1321
      10'd750  : in_data <= 14'h118f; // 'd4495
      10'd751  : in_data <= 14'h0a75; // 'd2677
      10'd752  : in_data <= 14'h0b08; // 'd2824
      10'd753  : in_data <= 14'h0356; // 'd854
      10'd754  : in_data <= 14'h0e64; // 'd3684
      10'd755  : in_data <= 14'h11d0; // 'd4560
      10'd756  : in_data <= 14'h0b43; // 'd2883
      10'd757  : in_data <= 14'h0889; // 'd2185
      10'd758  : in_data <= 14'h0462; // 'd1122
      10'd759  : in_data <= 14'h039a; // 'd922
      10'd760  : in_data <= 14'h12cf; // 'd4815
      10'd761  : in_data <= 14'h0b36; // 'd2870
      10'd762  : in_data <= 14'h0f6a; // 'd3946
      10'd763  : in_data <= 14'h0d7a; // 'd3450
      10'd764  : in_data <= 14'h07ed; // 'd2029
      10'd765  : in_data <= 14'h0084; // 'd132
      10'd766  : in_data <= 14'h037d; // 'd893
      10'd767  : in_data <= 14'h1384; // 'd4996
      10'd768  : in_data <= 14'h0cfa; // 'd3322
      10'd769  : in_data <= 14'h0ad6; // 'd2774
      10'd770  : in_data <= 14'h1301; // 'd4865
      10'd771  : in_data <= 14'h0762; // 'd1890
      10'd772  : in_data <= 14'h1126; // 'd4390
      10'd773  : in_data <= 14'h1213; // 'd4627
      10'd774  : in_data <= 14'h08f0; // 'd2288
      10'd775  : in_data <= 14'h0a5c; // 'd2652
      10'd776  : in_data <= 14'h007e; // 'd126
      10'd777  : in_data <= 14'h0acf; // 'd2767
      10'd778  : in_data <= 14'h0c15; // 'd3093
      10'd779  : in_data <= 14'h0898; // 'd2200
      10'd780  : in_data <= 14'h063a; // 'd1594
      10'd781  : in_data <= 14'h01d0; // 'd464
      10'd782  : in_data <= 14'h0954; // 'd2388
      10'd783  : in_data <= 14'h0789; // 'd1929
      10'd784  : in_data <= 14'h02aa; // 'd682
      10'd785  : in_data <= 14'h0858; // 'd2136
      10'd786  : in_data <= 14'h0962; // 'd2402
      10'd787  : in_data <= 14'h075d; // 'd1885
      10'd788  : in_data <= 14'h0be9; // 'd3049
      10'd789  : in_data <= 14'h01db; // 'd475
      10'd790  : in_data <= 14'h0dcf; // 'd3535
      10'd791  : in_data <= 14'h0245; // 'd581
      10'd792  : in_data <= 14'h0b3a; // 'd2874
      10'd793  : in_data <= 14'h03c6; // 'd966
      10'd794  : in_data <= 14'h092f; // 'd2351
      10'd795  : in_data <= 14'h06bb; // 'd1723
      10'd796  : in_data <= 14'h0590; // 'd1424
      10'd797  : in_data <= 14'h06ee; // 'd1774
      10'd798  : in_data <= 14'h00dc; // 'd220
      10'd799  : in_data <= 14'h0914; // 'd2324
      10'd800  : in_data <= 14'h005f; // 'd95
      10'd801  : in_data <= 14'h0aee; // 'd2798
      10'd802  : in_data <= 14'h03e3; // 'd995
      10'd803  : in_data <= 14'h0d30; // 'd3376
      10'd804  : in_data <= 14'h071c; // 'd1820
      10'd805  : in_data <= 14'h0e74; // 'd3700
      10'd806  : in_data <= 14'h0ac2; // 'd2754
      10'd807  : in_data <= 14'h0076; // 'd118
      10'd808  : in_data <= 14'h0954; // 'd2388
      10'd809  : in_data <= 14'h02b4; // 'd692
      10'd810  : in_data <= 14'h13cb; // 'd5067
      10'd811  : in_data <= 14'h115b; // 'd4443
      10'd812  : in_data <= 14'h13c9; // 'd5065
      10'd813  : in_data <= 14'h0d68; // 'd3432
      10'd814  : in_data <= 14'h002c; // 'd44
      10'd815  : in_data <= 14'h0056; // 'd86
      10'd816  : in_data <= 14'h05b4; // 'd1460
      10'd817  : in_data <= 14'h067a; // 'd1658
      10'd818  : in_data <= 14'h1137; // 'd4407
      10'd819  : in_data <= 14'h0f13; // 'd3859
      10'd820  : in_data <= 14'h10b2; // 'd4274
      10'd821  : in_data <= 14'h082e; // 'd2094
      10'd822  : in_data <= 14'h1330; // 'd4912
      10'd823  : in_data <= 14'h086f; // 'd2159
      10'd824  : in_data <= 14'h0979; // 'd2425
      10'd825  : in_data <= 14'h0d81; // 'd3457
      10'd826  : in_data <= 14'h0e5f; // 'd3679
      10'd827  : in_data <= 14'h10ac; // 'd4268
      10'd828  : in_data <= 14'h02cd; // 'd717
      10'd829  : in_data <= 14'h0d45; // 'd3397
      10'd830  : in_data <= 14'h1238; // 'd4664
      10'd831  : in_data <= 14'h11eb; // 'd4587
      10'd832  : in_data <= 14'h017d; // 'd381
      10'd833  : in_data <= 14'h006b; // 'd107
      10'd834  : in_data <= 14'h112a; // 'd4394
      10'd835  : in_data <= 14'h13f7; // 'd5111
      10'd836  : in_data <= 14'h0e35; // 'd3637
      10'd837  : in_data <= 14'h000e; // 'd14
      10'd838  : in_data <= 14'h0069; // 'd105
      10'd839  : in_data <= 14'h0124; // 'd292
      10'd840  : in_data <= 14'h004b; // 'd75
      10'd841  : in_data <= 14'h05c7; // 'd1479
      10'd842  : in_data <= 14'h1363; // 'd4963
      10'd843  : in_data <= 14'h11a9; // 'd4521
      10'd844  : in_data <= 14'h06a1; // 'd1697
      10'd845  : in_data <= 14'h069d; // 'd1693
      10'd846  : in_data <= 14'h1153; // 'd4435
      10'd847  : in_data <= 14'h04e1; // 'd1249
      10'd848  : in_data <= 14'h127b; // 'd4731
      10'd849  : in_data <= 14'h01c7; // 'd455
      10'd850  : in_data <= 14'h068e; // 'd1678
      10'd851  : in_data <= 14'h068b; // 'd1675
      10'd852  : in_data <= 14'h022f; // 'd559
      10'd853  : in_data <= 14'h0828; // 'd2088
      10'd854  : in_data <= 14'h08c7; // 'd2247
      10'd855  : in_data <= 14'h12bd; // 'd4797
      10'd856  : in_data <= 14'h0d7c; // 'd3452
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      11'd0    : out_data_ref <= 8'hf4;
      11'd1    : out_data_ref <= 8'h78;
      11'd2    : out_data_ref <= 8'h10;
      11'd3    : out_data_ref <= 8'h59;
      11'd4    : out_data_ref <= 8'he8;
      11'd5    : out_data_ref <= 8'h1a;
      11'd6    : out_data_ref <= 8'h38;
      11'd7    : out_data_ref <= 8'he6;
      11'd8    : out_data_ref <= 8'h78;
      11'd9    : out_data_ref <= 8'h9f;
      11'd10   : out_data_ref <= 8'h2f;
      11'd11   : out_data_ref <= 8'hc3;
      11'd12   : out_data_ref <= 8'h39;
      11'd13   : out_data_ref <= 8'h12;
      11'd14   : out_data_ref <= 8'he5;
      11'd15   : out_data_ref <= 8'h68;
      11'd16   : out_data_ref <= 8'hb5;
      11'd17   : out_data_ref <= 8'hb5;
      11'd18   : out_data_ref <= 8'he5;
      11'd19   : out_data_ref <= 8'hc5;
      11'd20   : out_data_ref <= 8'hc1;
      11'd21   : out_data_ref <= 8'hb0;
      11'd22   : out_data_ref <= 8'h4f;
      11'd23   : out_data_ref <= 8'h43;
      11'd24   : out_data_ref <= 8'hb6;
      11'd25   : out_data_ref <= 8'hde;
      11'd26   : out_data_ref <= 8'hd8;
      11'd27   : out_data_ref <= 8'h6a;
      11'd28   : out_data_ref <= 8'hc1;
      11'd29   : out_data_ref <= 8'hab;
      11'd30   : out_data_ref <= 8'hd4;
      11'd31   : out_data_ref <= 8'h30;
      11'd32   : out_data_ref <= 8'h47;
      11'd33   : out_data_ref <= 8'he5;
      11'd34   : out_data_ref <= 8'h55;
      11'd35   : out_data_ref <= 8'h37;
      11'd36   : out_data_ref <= 8'h0f;
      11'd37   : out_data_ref <= 8'hc9;
      11'd38   : out_data_ref <= 8'h57;
      11'd39   : out_data_ref <= 8'h96;
      11'd40   : out_data_ref <= 8'hae;
      11'd41   : out_data_ref <= 8'he8;
      11'd42   : out_data_ref <= 8'hc2;
      11'd43   : out_data_ref <= 8'hca;
      11'd44   : out_data_ref <= 8'h83;
      11'd45   : out_data_ref <= 8'hf1;
      11'd46   : out_data_ref <= 8'hd4;
      11'd47   : out_data_ref <= 8'h09;
      11'd48   : out_data_ref <= 8'h37;
      11'd49   : out_data_ref <= 8'h8e;
      11'd50   : out_data_ref <= 8'h23;
      11'd51   : out_data_ref <= 8'hf3;
      11'd52   : out_data_ref <= 8'ha9;
      11'd53   : out_data_ref <= 8'he7;
      11'd54   : out_data_ref <= 8'h75;
      11'd55   : out_data_ref <= 8'h95;
      11'd56   : out_data_ref <= 8'h85;
      11'd57   : out_data_ref <= 8'h6c;
      11'd58   : out_data_ref <= 8'h94;
      11'd59   : out_data_ref <= 8'hd9;
      11'd60   : out_data_ref <= 8'h56;
      11'd61   : out_data_ref <= 8'h34;
      11'd62   : out_data_ref <= 8'h6d;
      11'd63   : out_data_ref <= 8'h52;
      11'd64   : out_data_ref <= 8'h5a;
      11'd65   : out_data_ref <= 8'hf0;
      11'd66   : out_data_ref <= 8'h60;
      11'd67   : out_data_ref <= 8'h4e;
      11'd68   : out_data_ref <= 8'h5d;
      11'd69   : out_data_ref <= 8'hd1;
      11'd70   : out_data_ref <= 8'h6c;
      11'd71   : out_data_ref <= 8'h06;
      11'd72   : out_data_ref <= 8'h78;
      11'd73   : out_data_ref <= 8'hd6;
      11'd74   : out_data_ref <= 8'h7e;
      11'd75   : out_data_ref <= 8'h51;
      11'd76   : out_data_ref <= 8'h44;
      11'd77   : out_data_ref <= 8'h3c;
      11'd78   : out_data_ref <= 8'h60;
      11'd79   : out_data_ref <= 8'ha0;
      11'd80   : out_data_ref <= 8'hbb;
      11'd81   : out_data_ref <= 8'h21;
      11'd82   : out_data_ref <= 8'h99;
      11'd83   : out_data_ref <= 8'h39;
      11'd84   : out_data_ref <= 8'h4f;
      11'd85   : out_data_ref <= 8'h55;
      11'd86   : out_data_ref <= 8'ha8;
      11'd87   : out_data_ref <= 8'h1a;
      11'd88   : out_data_ref <= 8'h67;
      11'd89   : out_data_ref <= 8'h27;
      11'd90   : out_data_ref <= 8'h90;
      11'd91   : out_data_ref <= 8'h66;
      11'd92   : out_data_ref <= 8'hc4;
      11'd93   : out_data_ref <= 8'hf8;
      11'd94   : out_data_ref <= 8'h55;
      11'd95   : out_data_ref <= 8'h24;
      11'd96   : out_data_ref <= 8'h96;
      11'd97   : out_data_ref <= 8'h2a;
      11'd98   : out_data_ref <= 8'h78;
      11'd99   : out_data_ref <= 8'haf;
      11'd100  : out_data_ref <= 8'h51;
      11'd101  : out_data_ref <= 8'hb8;
      11'd102  : out_data_ref <= 8'h2e;
      11'd103  : out_data_ref <= 8'h2b;
      11'd104  : out_data_ref <= 8'h33;
      11'd105  : out_data_ref <= 8'hd7;
      11'd106  : out_data_ref <= 8'he8;
      11'd107  : out_data_ref <= 8'hb2;
      11'd108  : out_data_ref <= 8'h0d;
      11'd109  : out_data_ref <= 8'h0c;
      11'd110  : out_data_ref <= 8'hce;
      11'd111  : out_data_ref <= 8'h16;
      11'd112  : out_data_ref <= 8'hc2;
      11'd113  : out_data_ref <= 8'h3f;
      11'd114  : out_data_ref <= 8'h12;
      11'd115  : out_data_ref <= 8'h54;
      11'd116  : out_data_ref <= 8'hc9;
      11'd117  : out_data_ref <= 8'h20;
      11'd118  : out_data_ref <= 8'h25;
      11'd119  : out_data_ref <= 8'h2d;
      11'd120  : out_data_ref <= 8'he9;
      11'd121  : out_data_ref <= 8'h63;
      11'd122  : out_data_ref <= 8'h5e;
      11'd123  : out_data_ref <= 8'h3d;
      11'd124  : out_data_ref <= 8'h5d;
      11'd125  : out_data_ref <= 8'hb0;
      11'd126  : out_data_ref <= 8'h12;
      11'd127  : out_data_ref <= 8'h71;
      11'd128  : out_data_ref <= 8'h4d;
      11'd129  : out_data_ref <= 8'he3;
      11'd130  : out_data_ref <= 8'h4d;
      11'd131  : out_data_ref <= 8'h68;
      11'd132  : out_data_ref <= 8'hf4;
      11'd133  : out_data_ref <= 8'h33;
      11'd134  : out_data_ref <= 8'h34;
      11'd135  : out_data_ref <= 8'hf2;
      11'd136  : out_data_ref <= 8'hae;
      11'd137  : out_data_ref <= 8'ha8;
      11'd138  : out_data_ref <= 8'h0c;
      11'd139  : out_data_ref <= 8'h07;
      11'd140  : out_data_ref <= 8'hd2;
      11'd141  : out_data_ref <= 8'h6c;
      11'd142  : out_data_ref <= 8'hb7;
      11'd143  : out_data_ref <= 8'h82;
      11'd144  : out_data_ref <= 8'h29;
      11'd145  : out_data_ref <= 8'hb5;
      11'd146  : out_data_ref <= 8'ha0;
      11'd147  : out_data_ref <= 8'h04;
      11'd148  : out_data_ref <= 8'h0a;
      11'd149  : out_data_ref <= 8'h7c;
      11'd150  : out_data_ref <= 8'h44;
      11'd151  : out_data_ref <= 8'hfc;
      11'd152  : out_data_ref <= 8'h52;
      11'd153  : out_data_ref <= 8'h85;
      11'd154  : out_data_ref <= 8'hbd;
      11'd155  : out_data_ref <= 8'hd0;
      11'd156  : out_data_ref <= 8'h34;
      11'd157  : out_data_ref <= 8'h8c;
      11'd158  : out_data_ref <= 8'hb3;
      11'd159  : out_data_ref <= 8'h8f;
      11'd160  : out_data_ref <= 8'hcd;
      11'd161  : out_data_ref <= 8'h3b;
      11'd162  : out_data_ref <= 8'h84;
      11'd163  : out_data_ref <= 8'hdd;
      11'd164  : out_data_ref <= 8'h37;
      11'd165  : out_data_ref <= 8'h08;
      11'd166  : out_data_ref <= 8'hbe;
      11'd167  : out_data_ref <= 8'h88;
      11'd168  : out_data_ref <= 8'h43;
      11'd169  : out_data_ref <= 8'h9f;
      11'd170  : out_data_ref <= 8'h1f;
      11'd171  : out_data_ref <= 8'h92;
      11'd172  : out_data_ref <= 8'h8f;
      11'd173  : out_data_ref <= 8'h81;
      11'd174  : out_data_ref <= 8'h8d;
      11'd175  : out_data_ref <= 8'hf3;
      11'd176  : out_data_ref <= 8'hca;
      11'd177  : out_data_ref <= 8'h82;
      11'd178  : out_data_ref <= 8'hfb;
      11'd179  : out_data_ref <= 8'h50;
      11'd180  : out_data_ref <= 8'h3a;
      11'd181  : out_data_ref <= 8'h59;
      11'd182  : out_data_ref <= 8'h66;
      11'd183  : out_data_ref <= 8'h15;
      11'd184  : out_data_ref <= 8'he8;
      11'd185  : out_data_ref <= 8'h9d;
      11'd186  : out_data_ref <= 8'h1a;
      11'd187  : out_data_ref <= 8'h45;
      11'd188  : out_data_ref <= 8'hbd;
      11'd189  : out_data_ref <= 8'h4b;
      11'd190  : out_data_ref <= 8'hc4;
      11'd191  : out_data_ref <= 8'h1d;
      11'd192  : out_data_ref <= 8'hc0;
      11'd193  : out_data_ref <= 8'hdf;
      11'd194  : out_data_ref <= 8'hc3;
      11'd195  : out_data_ref <= 8'h84;
      11'd196  : out_data_ref <= 8'hf3;
      11'd197  : out_data_ref <= 8'hbc;
      11'd198  : out_data_ref <= 8'hf3;
      11'd199  : out_data_ref <= 8'h19;
      11'd200  : out_data_ref <= 8'h88;
      11'd201  : out_data_ref <= 8'h0a;
      11'd202  : out_data_ref <= 8'hf6;
      11'd203  : out_data_ref <= 8'h7f;
      11'd204  : out_data_ref <= 8'h4f;
      11'd205  : out_data_ref <= 8'h28;
      11'd206  : out_data_ref <= 8'h67;
      11'd207  : out_data_ref <= 8'h5e;
      11'd208  : out_data_ref <= 8'h58;
      11'd209  : out_data_ref <= 8'he2;
      11'd210  : out_data_ref <= 8'hbc;
      11'd211  : out_data_ref <= 8'h6a;
      11'd212  : out_data_ref <= 8'h85;
      11'd213  : out_data_ref <= 8'h89;
      11'd214  : out_data_ref <= 8'h1b;
      11'd215  : out_data_ref <= 8'hd3;
      11'd216  : out_data_ref <= 8'hd2;
      11'd217  : out_data_ref <= 8'h34;
      11'd218  : out_data_ref <= 8'hb7;
      11'd219  : out_data_ref <= 8'hc3;
      11'd220  : out_data_ref <= 8'h85;
      11'd221  : out_data_ref <= 8'hdd;
      11'd222  : out_data_ref <= 8'hb8;
      11'd223  : out_data_ref <= 8'h41;
      11'd224  : out_data_ref <= 8'h3a;
      11'd225  : out_data_ref <= 8'h0c;
      11'd226  : out_data_ref <= 8'hab;
      11'd227  : out_data_ref <= 8'h6d;
      11'd228  : out_data_ref <= 8'h20;
      11'd229  : out_data_ref <= 8'h85;
      11'd230  : out_data_ref <= 8'hb5;
      11'd231  : out_data_ref <= 8'h48;
      11'd232  : out_data_ref <= 8'hb0;
      11'd233  : out_data_ref <= 8'h7f;
      11'd234  : out_data_ref <= 8'h55;
      11'd235  : out_data_ref <= 8'hc9;
      11'd236  : out_data_ref <= 8'h08;
      11'd237  : out_data_ref <= 8'h21;
      11'd238  : out_data_ref <= 8'hf1;
      11'd239  : out_data_ref <= 8'hd3;
      11'd240  : out_data_ref <= 8'hd5;
      11'd241  : out_data_ref <= 8'h7d;
      11'd242  : out_data_ref <= 8'h5b;
      11'd243  : out_data_ref <= 8'h82;
      11'd244  : out_data_ref <= 8'h3b;
      11'd245  : out_data_ref <= 8'h54;
      11'd246  : out_data_ref <= 8'hd0;
      11'd247  : out_data_ref <= 8'h72;
      11'd248  : out_data_ref <= 8'h15;
      11'd249  : out_data_ref <= 8'h13;
      11'd250  : out_data_ref <= 8'h26;
      11'd251  : out_data_ref <= 8'h83;
      11'd252  : out_data_ref <= 8'h31;
      11'd253  : out_data_ref <= 8'hbe;
      11'd254  : out_data_ref <= 8'h37;
      11'd255  : out_data_ref <= 8'h14;
      11'd256  : out_data_ref <= 8'hc4;
      11'd257  : out_data_ref <= 8'heb;
      11'd258  : out_data_ref <= 8'h37;
      11'd259  : out_data_ref <= 8'h1c;
      11'd260  : out_data_ref <= 8'hbf;
      11'd261  : out_data_ref <= 8'h79;
      11'd262  : out_data_ref <= 8'h30;
      11'd263  : out_data_ref <= 8'h58;
      11'd264  : out_data_ref <= 8'h8f;
      11'd265  : out_data_ref <= 8'h5c;
      11'd266  : out_data_ref <= 8'h13;
      11'd267  : out_data_ref <= 8'h97;
      11'd268  : out_data_ref <= 8'h02;
      11'd269  : out_data_ref <= 8'h54;
      11'd270  : out_data_ref <= 8'hb5;
      11'd271  : out_data_ref <= 8'h70;
      11'd272  : out_data_ref <= 8'h26;
      11'd273  : out_data_ref <= 8'hd6;
      11'd274  : out_data_ref <= 8'h9a;
      11'd275  : out_data_ref <= 8'h56;
      11'd276  : out_data_ref <= 8'h84;
      11'd277  : out_data_ref <= 8'h09;
      11'd278  : out_data_ref <= 8'h02;
      11'd279  : out_data_ref <= 8'hf5;
      11'd280  : out_data_ref <= 8'h4e;
      11'd281  : out_data_ref <= 8'h7e;
      11'd282  : out_data_ref <= 8'hb6;
      11'd283  : out_data_ref <= 8'hc0;
      11'd284  : out_data_ref <= 8'hb5;
      11'd285  : out_data_ref <= 8'hfc;
      11'd286  : out_data_ref <= 8'hee;
      11'd287  : out_data_ref <= 8'hf1;
      11'd288  : out_data_ref <= 8'h82;
      11'd289  : out_data_ref <= 8'ha9;
      11'd290  : out_data_ref <= 8'h4b;
      11'd291  : out_data_ref <= 8'hff;
      11'd292  : out_data_ref <= 8'h67;
      11'd293  : out_data_ref <= 8'hd6;
      11'd294  : out_data_ref <= 8'ha0;
      11'd295  : out_data_ref <= 8'h9d;
      11'd296  : out_data_ref <= 8'h87;
      11'd297  : out_data_ref <= 8'hd7;
      11'd298  : out_data_ref <= 8'h2c;
      11'd299  : out_data_ref <= 8'hee;
      11'd300  : out_data_ref <= 8'h21;
      11'd301  : out_data_ref <= 8'h0f;
      11'd302  : out_data_ref <= 8'hd0;
      11'd303  : out_data_ref <= 8'h5b;
      11'd304  : out_data_ref <= 8'h69;
      11'd305  : out_data_ref <= 8'h66;
      11'd306  : out_data_ref <= 8'h5b;
      11'd307  : out_data_ref <= 8'he0;
      11'd308  : out_data_ref <= 8'he6;
      11'd309  : out_data_ref <= 8'had;
      11'd310  : out_data_ref <= 8'h1a;
      11'd311  : out_data_ref <= 8'hef;
      11'd312  : out_data_ref <= 8'heb;
      11'd313  : out_data_ref <= 8'hb5;
      11'd314  : out_data_ref <= 8'hc3;
      11'd315  : out_data_ref <= 8'hb5;
      11'd316  : out_data_ref <= 8'h29;
      11'd317  : out_data_ref <= 8'ha8;
      11'd318  : out_data_ref <= 8'h89;
      11'd319  : out_data_ref <= 8'hd3;
      11'd320  : out_data_ref <= 8'hcf;
      11'd321  : out_data_ref <= 8'h9e;
      11'd322  : out_data_ref <= 8'hfa;
      11'd323  : out_data_ref <= 8'ha3;
      11'd324  : out_data_ref <= 8'h8f;
      11'd325  : out_data_ref <= 8'h9b;
      11'd326  : out_data_ref <= 8'ha1;
      11'd327  : out_data_ref <= 8'h0a;
      11'd328  : out_data_ref <= 8'h97;
      11'd329  : out_data_ref <= 8'hfe;
      11'd330  : out_data_ref <= 8'hc6;
      11'd331  : out_data_ref <= 8'h87;
      11'd332  : out_data_ref <= 8'h43;
      11'd333  : out_data_ref <= 8'h07;
      11'd334  : out_data_ref <= 8'h53;
      11'd335  : out_data_ref <= 8'h13;
      11'd336  : out_data_ref <= 8'hd1;
      11'd337  : out_data_ref <= 8'h89;
      11'd338  : out_data_ref <= 8'h56;
      11'd339  : out_data_ref <= 8'h19;
      11'd340  : out_data_ref <= 8'h88;
      11'd341  : out_data_ref <= 8'h1a;
      11'd342  : out_data_ref <= 8'h77;
      11'd343  : out_data_ref <= 8'h6c;
      11'd344  : out_data_ref <= 8'he3;
      11'd345  : out_data_ref <= 8'h86;
      11'd346  : out_data_ref <= 8'hda;
      11'd347  : out_data_ref <= 8'hf1;
      11'd348  : out_data_ref <= 8'hd1;
      11'd349  : out_data_ref <= 8'h19;
      11'd350  : out_data_ref <= 8'h0c;
      11'd351  : out_data_ref <= 8'hfd;
      11'd352  : out_data_ref <= 8'h63;
      11'd353  : out_data_ref <= 8'h3f;
      11'd354  : out_data_ref <= 8'h88;
      11'd355  : out_data_ref <= 8'h70;
      11'd356  : out_data_ref <= 8'h3f;
      11'd357  : out_data_ref <= 8'h7e;
      11'd358  : out_data_ref <= 8'h42;
      11'd359  : out_data_ref <= 8'ha8;
      11'd360  : out_data_ref <= 8'h9a;
      11'd361  : out_data_ref <= 8'h07;
      11'd362  : out_data_ref <= 8'h92;
      11'd363  : out_data_ref <= 8'h35;
      11'd364  : out_data_ref <= 8'h01;
      11'd365  : out_data_ref <= 8'h28;
      11'd366  : out_data_ref <= 8'h86;
      11'd367  : out_data_ref <= 8'hfc;
      11'd368  : out_data_ref <= 8'hf1;
      11'd369  : out_data_ref <= 8'hc5;
      11'd370  : out_data_ref <= 8'hc6;
      11'd371  : out_data_ref <= 8'haa;
      11'd372  : out_data_ref <= 8'had;
      11'd373  : out_data_ref <= 8'h40;
      11'd374  : out_data_ref <= 8'h5f;
      11'd375  : out_data_ref <= 8'h6a;
      11'd376  : out_data_ref <= 8'hc3;
      11'd377  : out_data_ref <= 8'h80;
      11'd378  : out_data_ref <= 8'h39;
      11'd379  : out_data_ref <= 8'h2b;
      11'd380  : out_data_ref <= 8'h23;
      11'd381  : out_data_ref <= 8'h1e;
      11'd382  : out_data_ref <= 8'hb3;
      11'd383  : out_data_ref <= 8'hf8;
      11'd384  : out_data_ref <= 8'h16;
      11'd385  : out_data_ref <= 8'h3b;
      11'd386  : out_data_ref <= 8'haa;
      11'd387  : out_data_ref <= 8'he5;
      11'd388  : out_data_ref <= 8'h36;
      11'd389  : out_data_ref <= 8'hb9;
      11'd390  : out_data_ref <= 8'hbc;
      11'd391  : out_data_ref <= 8'h9d;
      11'd392  : out_data_ref <= 8'he5;
      11'd393  : out_data_ref <= 8'h52;
      11'd394  : out_data_ref <= 8'hcc;
      11'd395  : out_data_ref <= 8'h8c;
      11'd396  : out_data_ref <= 8'h81;
      11'd397  : out_data_ref <= 8'h3d;
      11'd398  : out_data_ref <= 8'h20;
      11'd399  : out_data_ref <= 8'h6a;
      11'd400  : out_data_ref <= 8'h65;
      11'd401  : out_data_ref <= 8'h9f;
      11'd402  : out_data_ref <= 8'hd3;
      11'd403  : out_data_ref <= 8'h04;
      11'd404  : out_data_ref <= 8'hb2;
      11'd405  : out_data_ref <= 8'h17;
      11'd406  : out_data_ref <= 8'hcb;
      11'd407  : out_data_ref <= 8'ha6;
      11'd408  : out_data_ref <= 8'h53;
      11'd409  : out_data_ref <= 8'h77;
      11'd410  : out_data_ref <= 8'h2c;
      11'd411  : out_data_ref <= 8'h7e;
      11'd412  : out_data_ref <= 8'h48;
      11'd413  : out_data_ref <= 8'h4a;
      11'd414  : out_data_ref <= 8'hec;
      11'd415  : out_data_ref <= 8'h75;
      11'd416  : out_data_ref <= 8'h32;
      11'd417  : out_data_ref <= 8'h9f;
      11'd418  : out_data_ref <= 8'hf7;
      11'd419  : out_data_ref <= 8'h84;
      11'd420  : out_data_ref <= 8'h1a;
      11'd421  : out_data_ref <= 8'h1d;
      11'd422  : out_data_ref <= 8'h97;
      11'd423  : out_data_ref <= 8'ha0;
      11'd424  : out_data_ref <= 8'h72;
      11'd425  : out_data_ref <= 8'h1b;
      11'd426  : out_data_ref <= 8'h99;
      11'd427  : out_data_ref <= 8'h65;
      11'd428  : out_data_ref <= 8'h63;
      11'd429  : out_data_ref <= 8'h70;
      11'd430  : out_data_ref <= 8'h40;
      11'd431  : out_data_ref <= 8'hea;
      11'd432  : out_data_ref <= 8'h10;
      11'd433  : out_data_ref <= 8'hd9;
      11'd434  : out_data_ref <= 8'hf6;
      11'd435  : out_data_ref <= 8'h2d;
      11'd436  : out_data_ref <= 8'haf;
      11'd437  : out_data_ref <= 8'h55;
      11'd438  : out_data_ref <= 8'he1;
      11'd439  : out_data_ref <= 8'h30;
      11'd440  : out_data_ref <= 8'ha4;
      11'd441  : out_data_ref <= 8'h4d;
      11'd442  : out_data_ref <= 8'he2;
      11'd443  : out_data_ref <= 8'h96;
      11'd444  : out_data_ref <= 8'h81;
      11'd445  : out_data_ref <= 8'h03;
      11'd446  : out_data_ref <= 8'hc2;
      11'd447  : out_data_ref <= 8'h37;
      11'd448  : out_data_ref <= 8'h6d;
      11'd449  : out_data_ref <= 8'h0f;
      11'd450  : out_data_ref <= 8'h21;
      11'd451  : out_data_ref <= 8'h05;
      11'd452  : out_data_ref <= 8'h66;
      11'd453  : out_data_ref <= 8'hb5;
      11'd454  : out_data_ref <= 8'hdf;
      11'd455  : out_data_ref <= 8'h98;
      11'd456  : out_data_ref <= 8'h7d;
      11'd457  : out_data_ref <= 8'hc3;
      11'd458  : out_data_ref <= 8'h74;
      11'd459  : out_data_ref <= 8'h7a;
      11'd460  : out_data_ref <= 8'h7b;
      11'd461  : out_data_ref <= 8'hf1;
      11'd462  : out_data_ref <= 8'hf8;
      11'd463  : out_data_ref <= 8'h50;
      11'd464  : out_data_ref <= 8'haf;
      11'd465  : out_data_ref <= 8'h40;
      11'd466  : out_data_ref <= 8'hae;
      11'd467  : out_data_ref <= 8'h4c;
      11'd468  : out_data_ref <= 8'h12;
      11'd469  : out_data_ref <= 8'h95;
      11'd470  : out_data_ref <= 8'h6f;
      11'd471  : out_data_ref <= 8'hf1;
      11'd472  : out_data_ref <= 8'hb4;
      11'd473  : out_data_ref <= 8'ha2;
      11'd474  : out_data_ref <= 8'hfe;
      11'd475  : out_data_ref <= 8'hc4;
      11'd476  : out_data_ref <= 8'h51;
      11'd477  : out_data_ref <= 8'hdf;
      11'd478  : out_data_ref <= 8'hb1;
      11'd479  : out_data_ref <= 8'h7e;
      11'd480  : out_data_ref <= 8'hdd;
      11'd481  : out_data_ref <= 8'hfe;
      11'd482  : out_data_ref <= 8'h7f;
      11'd483  : out_data_ref <= 8'h9a;
      11'd484  : out_data_ref <= 8'h46;
      11'd485  : out_data_ref <= 8'h31;
      11'd486  : out_data_ref <= 8'h23;
      11'd487  : out_data_ref <= 8'ha6;
      11'd488  : out_data_ref <= 8'hba;
      11'd489  : out_data_ref <= 8'h5d;
      11'd490  : out_data_ref <= 8'h65;
      11'd491  : out_data_ref <= 8'h1d;
      11'd492  : out_data_ref <= 8'he8;
      11'd493  : out_data_ref <= 8'h1a;
      11'd494  : out_data_ref <= 8'h58;
      11'd495  : out_data_ref <= 8'hf5;
      11'd496  : out_data_ref <= 8'h13;
      11'd497  : out_data_ref <= 8'hc6;
      11'd498  : out_data_ref <= 8'hb2;
      11'd499  : out_data_ref <= 8'h8f;
      11'd500  : out_data_ref <= 8'h28;
      11'd501  : out_data_ref <= 8'h14;
      11'd502  : out_data_ref <= 8'h8b;
      11'd503  : out_data_ref <= 8'h7f;
      11'd504  : out_data_ref <= 8'h42;
      11'd505  : out_data_ref <= 8'ha4;
      11'd506  : out_data_ref <= 8'hd5;
      11'd507  : out_data_ref <= 8'hcf;
      11'd508  : out_data_ref <= 8'h3e;
      11'd509  : out_data_ref <= 8'h7a;
      11'd510  : out_data_ref <= 8'h6a;
      11'd511  : out_data_ref <= 8'h84;
      11'd512  : out_data_ref <= 8'hcd;
      11'd513  : out_data_ref <= 8'h3b;
      11'd514  : out_data_ref <= 8'hf9;
      11'd515  : out_data_ref <= 8'h59;
      11'd516  : out_data_ref <= 8'h29;
      11'd517  : out_data_ref <= 8'h76;
      11'd518  : out_data_ref <= 8'h1d;
      11'd519  : out_data_ref <= 8'hae;
      11'd520  : out_data_ref <= 8'he5;
      11'd521  : out_data_ref <= 8'ha3;
      11'd522  : out_data_ref <= 8'h8e;
      11'd523  : out_data_ref <= 8'h1e;
      11'd524  : out_data_ref <= 8'h9a;
      11'd525  : out_data_ref <= 8'hd0;
      11'd526  : out_data_ref <= 8'h6c;
      11'd527  : out_data_ref <= 8'h6a;
      11'd528  : out_data_ref <= 8'h69;
      11'd529  : out_data_ref <= 8'h32;
      11'd530  : out_data_ref <= 8'hbf;
      11'd531  : out_data_ref <= 8'h04;
      11'd532  : out_data_ref <= 8'he3;
      11'd533  : out_data_ref <= 8'h71;
      11'd534  : out_data_ref <= 8'hca;
      11'd535  : out_data_ref <= 8'hf5;
      11'd536  : out_data_ref <= 8'hc1;
      11'd537  : out_data_ref <= 8'h05;
      11'd538  : out_data_ref <= 8'h12;
      11'd539  : out_data_ref <= 8'h19;
      11'd540  : out_data_ref <= 8'h07;
      11'd541  : out_data_ref <= 8'h39;
      11'd542  : out_data_ref <= 8'hea;
      11'd543  : out_data_ref <= 8'h5a;
      11'd544  : out_data_ref <= 8'h90;
      11'd545  : out_data_ref <= 8'h62;
      11'd546  : out_data_ref <= 8'h55;
      11'd547  : out_data_ref <= 8'h8b;
      11'd548  : out_data_ref <= 8'hc0;
      11'd549  : out_data_ref <= 8'h50;
      11'd550  : out_data_ref <= 8'ha0;
      11'd551  : out_data_ref <= 8'hdd;
      11'd552  : out_data_ref <= 8'h2a;
      11'd553  : out_data_ref <= 8'hf1;
      11'd554  : out_data_ref <= 8'h73;
      11'd555  : out_data_ref <= 8'h75;
      11'd556  : out_data_ref <= 8'h69;
      11'd557  : out_data_ref <= 8'h1a;
      11'd558  : out_data_ref <= 8'h70;
      11'd559  : out_data_ref <= 8'h74;
      11'd560  : out_data_ref <= 8'h3d;
      11'd561  : out_data_ref <= 8'he9;
      11'd562  : out_data_ref <= 8'h25;
      11'd563  : out_data_ref <= 8'h4c;
      11'd564  : out_data_ref <= 8'hc5;
      11'd565  : out_data_ref <= 8'h40;
      11'd566  : out_data_ref <= 8'he1;
      11'd567  : out_data_ref <= 8'h15;
      11'd568  : out_data_ref <= 8'ha9;
      11'd569  : out_data_ref <= 8'h6f;
      11'd570  : out_data_ref <= 8'hb5;
      11'd571  : out_data_ref <= 8'h7c;
      11'd572  : out_data_ref <= 8'h27;
      11'd573  : out_data_ref <= 8'h58;
      11'd574  : out_data_ref <= 8'h8f;
      11'd575  : out_data_ref <= 8'hac;
      11'd576  : out_data_ref <= 8'h56;
      11'd577  : out_data_ref <= 8'hc9;
      11'd578  : out_data_ref <= 8'hfd;
      11'd579  : out_data_ref <= 8'he9;
      11'd580  : out_data_ref <= 8'he9;
      11'd581  : out_data_ref <= 8'h32;
      11'd582  : out_data_ref <= 8'h45;
      11'd583  : out_data_ref <= 8'hcc;
      11'd584  : out_data_ref <= 8'hae;
      11'd585  : out_data_ref <= 8'hce;
      11'd586  : out_data_ref <= 8'ha1;
      11'd587  : out_data_ref <= 8'hd1;
      11'd588  : out_data_ref <= 8'h0d;
      11'd589  : out_data_ref <= 8'h73;
      11'd590  : out_data_ref <= 8'hda;
      11'd591  : out_data_ref <= 8'h47;
      11'd592  : out_data_ref <= 8'h1f;
      11'd593  : out_data_ref <= 8'h28;
      11'd594  : out_data_ref <= 8'h05;
      11'd595  : out_data_ref <= 8'h5c;
      11'd596  : out_data_ref <= 8'h0f;
      11'd597  : out_data_ref <= 8'ha7;
      11'd598  : out_data_ref <= 8'hef;
      11'd599  : out_data_ref <= 8'h59;
      11'd600  : out_data_ref <= 8'h03;
      11'd601  : out_data_ref <= 8'hc5;
      11'd602  : out_data_ref <= 8'h91;
      11'd603  : out_data_ref <= 8'h5a;
      11'd604  : out_data_ref <= 8'hf1;
      11'd605  : out_data_ref <= 8'hc7;
      11'd606  : out_data_ref <= 8'h49;
      11'd607  : out_data_ref <= 8'h6f;
      11'd608  : out_data_ref <= 8'hd0;
      11'd609  : out_data_ref <= 8'hdf;
      11'd610  : out_data_ref <= 8'h17;
      11'd611  : out_data_ref <= 8'hcf;
      11'd612  : out_data_ref <= 8'h53;
      11'd613  : out_data_ref <= 8'h3a;
      11'd614  : out_data_ref <= 8'h48;
      11'd615  : out_data_ref <= 8'h0d;
      11'd616  : out_data_ref <= 8'h6b;
      11'd617  : out_data_ref <= 8'hde;
      11'd618  : out_data_ref <= 8'h7e;
      11'd619  : out_data_ref <= 8'hb2;
      11'd620  : out_data_ref <= 8'h91;
      11'd621  : out_data_ref <= 8'hd7;
      11'd622  : out_data_ref <= 8'h00;
      11'd623  : out_data_ref <= 8'h0d;
      11'd624  : out_data_ref <= 8'h74;
      11'd625  : out_data_ref <= 8'h70;
      11'd626  : out_data_ref <= 8'hca;
      11'd627  : out_data_ref <= 8'h0c;
      11'd628  : out_data_ref <= 8'h7d;
      11'd629  : out_data_ref <= 8'h35;
      11'd630  : out_data_ref <= 8'h0f;
      11'd631  : out_data_ref <= 8'hd1;
      11'd632  : out_data_ref <= 8'h75;
      11'd633  : out_data_ref <= 8'ha8;
      11'd634  : out_data_ref <= 8'hd4;
      11'd635  : out_data_ref <= 8'h6f;
      11'd636  : out_data_ref <= 8'hfc;
      11'd637  : out_data_ref <= 8'hfd;
      11'd638  : out_data_ref <= 8'h94;
      11'd639  : out_data_ref <= 8'h2a;
      11'd640  : out_data_ref <= 8'hf5;
      11'd641  : out_data_ref <= 8'h96;
      11'd642  : out_data_ref <= 8'h48;
      11'd643  : out_data_ref <= 8'h78;
      11'd644  : out_data_ref <= 8'hc5;
      11'd645  : out_data_ref <= 8'h60;
      11'd646  : out_data_ref <= 8'hd2;
      11'd647  : out_data_ref <= 8'h7c;
      11'd648  : out_data_ref <= 8'h44;
      11'd649  : out_data_ref <= 8'h92;
      11'd650  : out_data_ref <= 8'h07;
      11'd651  : out_data_ref <= 8'h7d;
      11'd652  : out_data_ref <= 8'hfa;
      11'd653  : out_data_ref <= 8'h0e;
      11'd654  : out_data_ref <= 8'hbb;
      11'd655  : out_data_ref <= 8'ha4;
      11'd656  : out_data_ref <= 8'h3d;
      11'd657  : out_data_ref <= 8'ha9;
      11'd658  : out_data_ref <= 8'hc7;
      11'd659  : out_data_ref <= 8'hde;
      11'd660  : out_data_ref <= 8'h44;
      11'd661  : out_data_ref <= 8'h1d;
      11'd662  : out_data_ref <= 8'hda;
      11'd663  : out_data_ref <= 8'h8a;
      11'd664  : out_data_ref <= 8'had;
      11'd665  : out_data_ref <= 8'ha7;
      11'd666  : out_data_ref <= 8'ha4;
      11'd667  : out_data_ref <= 8'h3b;
      11'd668  : out_data_ref <= 8'h93;
      11'd669  : out_data_ref <= 8'hf8;
      11'd670  : out_data_ref <= 8'h63;
      11'd671  : out_data_ref <= 8'h7d;
      11'd672  : out_data_ref <= 8'h79;
      11'd673  : out_data_ref <= 8'h8c;
      11'd674  : out_data_ref <= 8'h9b;
      11'd675  : out_data_ref <= 8'h5d;
      11'd676  : out_data_ref <= 8'h94;
      11'd677  : out_data_ref <= 8'h9e;
      11'd678  : out_data_ref <= 8'hf6;
      11'd679  : out_data_ref <= 8'h8c;
      11'd680  : out_data_ref <= 8'he1;
      11'd681  : out_data_ref <= 8'hda;
      11'd682  : out_data_ref <= 8'h51;
      11'd683  : out_data_ref <= 8'h36;
      11'd684  : out_data_ref <= 8'hfc;
      11'd685  : out_data_ref <= 8'h13;
      11'd686  : out_data_ref <= 8'hd6;
      11'd687  : out_data_ref <= 8'h54;
      11'd688  : out_data_ref <= 8'haf;
      11'd689  : out_data_ref <= 8'h82;
      11'd690  : out_data_ref <= 8'h0b;
      11'd691  : out_data_ref <= 8'hb1;
      11'd692  : out_data_ref <= 8'h62;
      11'd693  : out_data_ref <= 8'h0e;
      11'd694  : out_data_ref <= 8'hb5;
      11'd695  : out_data_ref <= 8'h35;
      11'd696  : out_data_ref <= 8'h87;
      11'd697  : out_data_ref <= 8'h81;
      11'd698  : out_data_ref <= 8'h04;
      11'd699  : out_data_ref <= 8'h69;
      11'd700  : out_data_ref <= 8'h4f;
      11'd701  : out_data_ref <= 8'h5a;
      11'd702  : out_data_ref <= 8'hd4;
      11'd703  : out_data_ref <= 8'h22;
      11'd704  : out_data_ref <= 8'ha4;
      11'd705  : out_data_ref <= 8'h8d;
      11'd706  : out_data_ref <= 8'h45;
      11'd707  : out_data_ref <= 8'h27;
      11'd708  : out_data_ref <= 8'he0;
      11'd709  : out_data_ref <= 8'hbb;
      11'd710  : out_data_ref <= 8'hd3;
      11'd711  : out_data_ref <= 8'h35;
      11'd712  : out_data_ref <= 8'h7d;
      11'd713  : out_data_ref <= 8'hac;
      11'd714  : out_data_ref <= 8'h6f;
      11'd715  : out_data_ref <= 8'h3f;
      11'd716  : out_data_ref <= 8'h43;
      11'd717  : out_data_ref <= 8'h3a;
      11'd718  : out_data_ref <= 8'h58;
      11'd719  : out_data_ref <= 8'hd0;
      11'd720  : out_data_ref <= 8'h65;
      11'd721  : out_data_ref <= 8'h2e;
      11'd722  : out_data_ref <= 8'h43;
      11'd723  : out_data_ref <= 8'h22;
      11'd724  : out_data_ref <= 8'heb;
      11'd725  : out_data_ref <= 8'hc3;
      11'd726  : out_data_ref <= 8'h46;
      11'd727  : out_data_ref <= 8'hfa;
      11'd728  : out_data_ref <= 8'h04;
      11'd729  : out_data_ref <= 8'h40;
      11'd730  : out_data_ref <= 8'hff;
      11'd731  : out_data_ref <= 8'h1f;
      11'd732  : out_data_ref <= 8'h62;
      11'd733  : out_data_ref <= 8'hec;
      11'd734  : out_data_ref <= 8'ha6;
      11'd735  : out_data_ref <= 8'h7a;
      11'd736  : out_data_ref <= 8'h8e;
      11'd737  : out_data_ref <= 8'h46;
      11'd738  : out_data_ref <= 8'hfd;
      11'd739  : out_data_ref <= 8'h96;
      11'd740  : out_data_ref <= 8'h09;
      11'd741  : out_data_ref <= 8'hcc;
      11'd742  : out_data_ref <= 8'hdc;
      11'd743  : out_data_ref <= 8'h66;
      11'd744  : out_data_ref <= 8'h5b;
      11'd745  : out_data_ref <= 8'h40;
      11'd746  : out_data_ref <= 8'hd6;
      11'd747  : out_data_ref <= 8'h40;
      11'd748  : out_data_ref <= 8'hcd;
      11'd749  : out_data_ref <= 8'h2b;
      11'd750  : out_data_ref <= 8'h0a;
      11'd751  : out_data_ref <= 8'h21;
      11'd752  : out_data_ref <= 8'hd2;
      11'd753  : out_data_ref <= 8'h5f;
      11'd754  : out_data_ref <= 8'h94;
      11'd755  : out_data_ref <= 8'h93;
      11'd756  : out_data_ref <= 8'h6a;
      11'd757  : out_data_ref <= 8'h50;
      11'd758  : out_data_ref <= 8'ha8;
      11'd759  : out_data_ref <= 8'hb5;
      11'd760  : out_data_ref <= 8'hb9;
      11'd761  : out_data_ref <= 8'h59;
      11'd762  : out_data_ref <= 8'hd0;
      11'd763  : out_data_ref <= 8'h10;
      11'd764  : out_data_ref <= 8'h29;
      11'd765  : out_data_ref <= 8'h70;
      11'd766  : out_data_ref <= 8'hb9;
      11'd767  : out_data_ref <= 8'he8;
      11'd768  : out_data_ref <= 8'h44;
      11'd769  : out_data_ref <= 8'hc2;
      11'd770  : out_data_ref <= 8'hff;
      11'd771  : out_data_ref <= 8'h15;
      11'd772  : out_data_ref <= 8'ha3;
      11'd773  : out_data_ref <= 8'hde;
      11'd774  : out_data_ref <= 8'hd4;
      11'd775  : out_data_ref <= 8'h1f;
      11'd776  : out_data_ref <= 8'h7f;
      11'd777  : out_data_ref <= 8'h28;
      11'd778  : out_data_ref <= 8'hfd;
      11'd779  : out_data_ref <= 8'h7f;
      11'd780  : out_data_ref <= 8'h6a;
      11'd781  : out_data_ref <= 8'h9b;
      11'd782  : out_data_ref <= 8'h7b;
      11'd783  : out_data_ref <= 8'h1f;
      11'd784  : out_data_ref <= 8'hd2;
      11'd785  : out_data_ref <= 8'h6a;
      11'd786  : out_data_ref <= 8'h75;
      11'd787  : out_data_ref <= 8'ha7;
      11'd788  : out_data_ref <= 8'h1e;
      11'd789  : out_data_ref <= 8'h7f;
      11'd790  : out_data_ref <= 8'h7a;
      11'd791  : out_data_ref <= 8'hdc;
      11'd792  : out_data_ref <= 8'h94;
      11'd793  : out_data_ref <= 8'h34;
      11'd794  : out_data_ref <= 8'h84;
      11'd795  : out_data_ref <= 8'he1;
      11'd796  : out_data_ref <= 8'h42;
      11'd797  : out_data_ref <= 8'he3;
      11'd798  : out_data_ref <= 8'h88;
      11'd799  : out_data_ref <= 8'h3b;
      11'd800  : out_data_ref <= 8'h11;
      11'd801  : out_data_ref <= 8'h9a;
      11'd802  : out_data_ref <= 8'hb3;
      11'd803  : out_data_ref <= 8'h2f;
      11'd804  : out_data_ref <= 8'h68;
      11'd805  : out_data_ref <= 8'hbe;
      11'd806  : out_data_ref <= 8'h6c;
      11'd807  : out_data_ref <= 8'h58;
      11'd808  : out_data_ref <= 8'h60;
      11'd809  : out_data_ref <= 8'h98;
      11'd810  : out_data_ref <= 8'h80;
      11'd811  : out_data_ref <= 8'h5f;
      11'd812  : out_data_ref <= 8'he1;
      11'd813  : out_data_ref <= 8'ha9;
      11'd814  : out_data_ref <= 8'hf6;
      11'd815  : out_data_ref <= 8'hc7;
      11'd816  : out_data_ref <= 8'h1a;
      11'd817  : out_data_ref <= 8'hbe;
      11'd818  : out_data_ref <= 8'hb4;
      11'd819  : out_data_ref <= 8'h51;
      11'd820  : out_data_ref <= 8'h24;
      11'd821  : out_data_ref <= 8'h29;
      11'd822  : out_data_ref <= 8'h91;
      11'd823  : out_data_ref <= 8'h4b;
      11'd824  : out_data_ref <= 8'h28;
      11'd825  : out_data_ref <= 8'h98;
      11'd826  : out_data_ref <= 8'hf3;
      11'd827  : out_data_ref <= 8'h8d;
      11'd828  : out_data_ref <= 8'h78;
      11'd829  : out_data_ref <= 8'hd6;
      11'd830  : out_data_ref <= 8'h5d;
      11'd831  : out_data_ref <= 8'hb8;
      11'd832  : out_data_ref <= 8'h22;
      11'd833  : out_data_ref <= 8'h71;
      11'd834  : out_data_ref <= 8'h83;
      11'd835  : out_data_ref <= 8'h07;
      11'd836  : out_data_ref <= 8'hc7;
      11'd837  : out_data_ref <= 8'h28;
      11'd838  : out_data_ref <= 8'h05;
      11'd839  : out_data_ref <= 8'h06;
      11'd840  : out_data_ref <= 8'hd4;
      11'd841  : out_data_ref <= 8'h9b;
      11'd842  : out_data_ref <= 8'h6a;
      11'd843  : out_data_ref <= 8'h85;
      11'd844  : out_data_ref <= 8'h74;
      11'd845  : out_data_ref <= 8'h81;
      11'd846  : out_data_ref <= 8'ha2;
      11'd847  : out_data_ref <= 8'h8a;
      11'd848  : out_data_ref <= 8'h04;
      11'd849  : out_data_ref <= 8'hf2;
      11'd850  : out_data_ref <= 8'h13;
      11'd851  : out_data_ref <= 8'h16;
      11'd852  : out_data_ref <= 8'h87;
      11'd853  : out_data_ref <= 8'ha1;
      11'd854  : out_data_ref <= 8'h7a;
      11'd855  : out_data_ref <= 8'h3d;
      11'd856  : out_data_ref <= 8'h04;
      11'd857  : out_data_ref <= 8'h63;
      11'd858  : out_data_ref <= 8'he3;
      11'd859  : out_data_ref <= 8'hcd;
      11'd860  : out_data_ref <= 8'h39;
      11'd861  : out_data_ref <= 8'h29;
      11'd862  : out_data_ref <= 8'hbc;
      11'd863  : out_data_ref <= 8'hbb;
      11'd864  : out_data_ref <= 8'h87;
      11'd865  : out_data_ref <= 8'h7b;
      11'd866  : out_data_ref <= 8'hbd;
      11'd867  : out_data_ref <= 8'hbc;
      11'd868  : out_data_ref <= 8'h52;
      11'd869  : out_data_ref <= 8'h60;
      11'd870  : out_data_ref <= 8'h6e;
      11'd871  : out_data_ref <= 8'h36;
      11'd872  : out_data_ref <= 8'h81;
      11'd873  : out_data_ref <= 8'h1e;
      11'd874  : out_data_ref <= 8'h96;
      11'd875  : out_data_ref <= 8'he6;
      11'd876  : out_data_ref <= 8'h9c;
      11'd877  : out_data_ref <= 8'he0;
      11'd878  : out_data_ref <= 8'hff;
      11'd879  : out_data_ref <= 8'h88;
      11'd880  : out_data_ref <= 8'h12;
      11'd881  : out_data_ref <= 8'hf3;
      11'd882  : out_data_ref <= 8'h0e;
      11'd883  : out_data_ref <= 8'h4a;
      11'd884  : out_data_ref <= 8'h6f;
      11'd885  : out_data_ref <= 8'h75;
      11'd886  : out_data_ref <= 8'h22;
      11'd887  : out_data_ref <= 8'he7;
      11'd888  : out_data_ref <= 8'h60;
      11'd889  : out_data_ref <= 8'h1e;
      11'd890  : out_data_ref <= 8'h31;
      11'd891  : out_data_ref <= 8'hf6;
      11'd892  : out_data_ref <= 8'h9e;
      11'd893  : out_data_ref <= 8'h3a;
      11'd894  : out_data_ref <= 8'h0b;
      11'd895  : out_data_ref <= 8'h8c;
      11'd896  : out_data_ref <= 8'hc3;
      11'd897  : out_data_ref <= 8'h00;
      11'd898  : out_data_ref <= 8'h0b;
      11'd899  : out_data_ref <= 8'hb3;
      11'd900  : out_data_ref <= 8'hce;
      11'd901  : out_data_ref <= 8'h5f;
      11'd902  : out_data_ref <= 8'h39;
      11'd903  : out_data_ref <= 8'hdd;
      11'd904  : out_data_ref <= 8'h47;
      11'd905  : out_data_ref <= 8'h7c;
      11'd906  : out_data_ref <= 8'hf0;
      11'd907  : out_data_ref <= 8'h28;
      11'd908  : out_data_ref <= 8'h97;
      11'd909  : out_data_ref <= 8'hd1;
      11'd910  : out_data_ref <= 8'h8d;
      11'd911  : out_data_ref <= 8'haa;
      11'd912  : out_data_ref <= 8'h2e;
      11'd913  : out_data_ref <= 8'hdf;
      11'd914  : out_data_ref <= 8'hec;
      11'd915  : out_data_ref <= 8'h88;
      11'd916  : out_data_ref <= 8'hdf;
      11'd917  : out_data_ref <= 8'h54;
      11'd918  : out_data_ref <= 8'h2a;
      11'd919  : out_data_ref <= 8'h8a;
      11'd920  : out_data_ref <= 8'h0c;
      11'd921  : out_data_ref <= 8'hb5;
      11'd922  : out_data_ref <= 8'he1;
      11'd923  : out_data_ref <= 8'h49;
      11'd924  : out_data_ref <= 8'h2e;
      11'd925  : out_data_ref <= 8'h48;
      11'd926  : out_data_ref <= 8'h6f;
      11'd927  : out_data_ref <= 8'h31;
      11'd928  : out_data_ref <= 8'h4d;
      11'd929  : out_data_ref <= 8'h88;
      11'd930  : out_data_ref <= 8'h9e;
      11'd931  : out_data_ref <= 8'h1d;
      11'd932  : out_data_ref <= 8'h2b;
      11'd933  : out_data_ref <= 8'hf6;
      11'd934  : out_data_ref <= 8'hba;
      11'd935  : out_data_ref <= 8'h8d;
      11'd936  : out_data_ref <= 8'ha3;
      11'd937  : out_data_ref <= 8'h50;
      11'd938  : out_data_ref <= 8'hf3;
      11'd939  : out_data_ref <= 8'hc0;
      11'd940  : out_data_ref <= 8'hb6;
      11'd941  : out_data_ref <= 8'hcb;
      11'd942  : out_data_ref <= 8'h32;
      11'd943  : out_data_ref <= 8'ha1;
      11'd944  : out_data_ref <= 8'h93;
      11'd945  : out_data_ref <= 8'h12;
      11'd946  : out_data_ref <= 8'hb3;
      11'd947  : out_data_ref <= 8'hbf;
      11'd948  : out_data_ref <= 8'h61;
      11'd949  : out_data_ref <= 8'h89;
      11'd950  : out_data_ref <= 8'h2e;
      11'd951  : out_data_ref <= 8'h54;
      11'd952  : out_data_ref <= 8'h6a;
      11'd953  : out_data_ref <= 8'h99;
      11'd954  : out_data_ref <= 8'h52;
      11'd955  : out_data_ref <= 8'h2f;
      11'd956  : out_data_ref <= 8'heb;
      11'd957  : out_data_ref <= 8'h4c;
      11'd958  : out_data_ref <= 8'hc8;
      11'd959  : out_data_ref <= 8'h5b;
      11'd960  : out_data_ref <= 8'h01;
      11'd961  : out_data_ref <= 8'h8c;
      11'd962  : out_data_ref <= 8'h8e;
      11'd963  : out_data_ref <= 8'h36;
      11'd964  : out_data_ref <= 8'he8;
      11'd965  : out_data_ref <= 8'h08;
      11'd966  : out_data_ref <= 8'h84;
      11'd967  : out_data_ref <= 8'h28;
      11'd968  : out_data_ref <= 8'h3b;
      11'd969  : out_data_ref <= 8'h1a;
      11'd970  : out_data_ref <= 8'h77;
      11'd971  : out_data_ref <= 8'h06;
      11'd972  : out_data_ref <= 8'h01;
      11'd973  : out_data_ref <= 8'h94;
      11'd974  : out_data_ref <= 8'h2d;
      11'd975  : out_data_ref <= 8'h50;
      11'd976  : out_data_ref <= 8'h60;
      11'd977  : out_data_ref <= 8'h1b;
      11'd978  : out_data_ref <= 8'h19;
      11'd979  : out_data_ref <= 8'ha0;
      11'd980  : out_data_ref <= 8'hac;
      11'd981  : out_data_ref <= 8'hb4;
      11'd982  : out_data_ref <= 8'h0e;
      11'd983  : out_data_ref <= 8'h44;
      11'd984  : out_data_ref <= 8'h90;
      11'd985  : out_data_ref <= 8'h70;
      11'd986  : out_data_ref <= 8'h48;
      11'd987  : out_data_ref <= 8'h8e;
      11'd988  : out_data_ref <= 8'haa;
      11'd989  : out_data_ref <= 8'h2d;
      11'd990  : out_data_ref <= 8'hb0;
      11'd991  : out_data_ref <= 8'h69;
      11'd992  : out_data_ref <= 8'hcf;
      11'd993  : out_data_ref <= 8'h2c;
      11'd994  : out_data_ref <= 8'hda;
      11'd995  : out_data_ref <= 8'h25;
      11'd996  : out_data_ref <= 8'h12;
      11'd997  : out_data_ref <= 8'h01;
      11'd998  : out_data_ref <= 8'had;
      11'd999  : out_data_ref <= 8'hda;
      11'd1000 : out_data_ref <= 8'hbe;
      11'd1001 : out_data_ref <= 8'hda;
      11'd1002 : out_data_ref <= 8'h2f;
      11'd1003 : out_data_ref <= 8'h84;
      11'd1004 : out_data_ref <= 8'h38;
      11'd1005 : out_data_ref <= 8'h16;
      11'd1006 : out_data_ref <= 8'h0f;
      11'd1007 : out_data_ref <= 8'h98;
      11'd1008 : out_data_ref <= 8'hf2;
      11'd1009 : out_data_ref <= 8'h40;
      11'd1010 : out_data_ref <= 8'h29;
      11'd1011 : out_data_ref <= 8'he4;
      11'd1012 : out_data_ref <= 8'hfe;
      11'd1013 : out_data_ref <= 8'he3;
      11'd1014 : out_data_ref <= 8'hea;
      11'd1015 : out_data_ref <= 8'h7f;
      11'd1016 : out_data_ref <= 8'hd1;
      11'd1017 : out_data_ref <= 8'h52;
      11'd1018 : out_data_ref <= 8'h6e;
      11'd1019 : out_data_ref <= 8'h5c;
      11'd1020 : out_data_ref <= 8'hbc;
      11'd1021 : out_data_ref <= 8'hde;
      11'd1022 : out_data_ref <= 8'h08;
      11'd1023 : out_data_ref <= 8'hc6;
      11'd1024 : out_data_ref <= 8'h99;
      11'd1025 : out_data_ref <= 8'h9f;
      11'd1026 : out_data_ref <= 8'h7e;
      11'd1027 : out_data_ref <= 8'h75;
      11'd1028 : out_data_ref <= 8'hc6;
      11'd1029 : out_data_ref <= 8'hb8;
      11'd1030 : out_data_ref <= 8'h7e;
      11'd1031 : out_data_ref <= 8'hf7;
      11'd1032 : out_data_ref <= 8'hf7;
      11'd1033 : out_data_ref <= 8'h3d;
      11'd1034 : out_data_ref <= 8'h6b;
      11'd1035 : out_data_ref <= 8'h87;
      11'd1036 : out_data_ref <= 8'h82;
      11'd1037 : out_data_ref <= 8'h1e;
      11'd1038 : out_data_ref <= 8'hd9;
      11'd1039 : out_data_ref <= 8'h20;
      11'd1040 : out_data_ref <= 8'h15;
      11'd1041 : out_data_ref <= 8'hd1;
      11'd1042 : out_data_ref <= 8'h6d;
      11'd1043 : out_data_ref <= 8'hb0;
      11'd1044 : out_data_ref <= 8'h6b;
      11'd1045 : out_data_ref <= 8'h6c;
      11'd1046 : out_data_ref <= 8'h62;
      11'd1047 : out_data_ref <= 8'h62;
      11'd1048 : out_data_ref <= 8'h52;
      11'd1049 : out_data_ref <= 8'h84;
      11'd1050 : out_data_ref <= 8'h92;
      11'd1051 : out_data_ref <= 8'h64;
      11'd1052 : out_data_ref <= 8'h88;
      11'd1053 : out_data_ref <= 8'hdd;
      11'd1054 : out_data_ref <= 8'h74;
      11'd1055 : out_data_ref <= 8'h33;
      11'd1056 : out_data_ref <= 8'hcc;
      11'd1057 : out_data_ref <= 8'h7b;
      11'd1058 : out_data_ref <= 8'h06;
      11'd1059 : out_data_ref <= 8'h9e;
      11'd1060 : out_data_ref <= 8'h02;
      11'd1061 : out_data_ref <= 8'h95;
      11'd1062 : out_data_ref <= 8'h90;
      11'd1063 : out_data_ref <= 8'h63;
      11'd1064 : out_data_ref <= 8'h50;
      11'd1065 : out_data_ref <= 8'ha9;
      11'd1066 : out_data_ref <= 8'hd4;
      11'd1067 : out_data_ref <= 8'hb5;
      11'd1068 : out_data_ref <= 8'h83;
      11'd1069 : out_data_ref <= 8'h14;
      11'd1070 : out_data_ref <= 8'h70;
      11'd1071 : out_data_ref <= 8'h9a;
      11'd1072 : out_data_ref <= 8'h09;
      11'd1073 : out_data_ref <= 8'hd9;
      11'd1074 : out_data_ref <= 8'h1b;
      11'd1075 : out_data_ref <= 8'hf6;
      11'd1076 : out_data_ref <= 8'h2a;
      11'd1077 : out_data_ref <= 8'h59;
      11'd1078 : out_data_ref <= 8'h82;
      11'd1079 : out_data_ref <= 8'h7d;
      11'd1080 : out_data_ref <= 8'h61;
      11'd1081 : out_data_ref <= 8'h97;
      11'd1082 : out_data_ref <= 8'hfd;
      11'd1083 : out_data_ref <= 8'h8d;
      11'd1084 : out_data_ref <= 8'h91;
      11'd1085 : out_data_ref <= 8'hb4;
      11'd1086 : out_data_ref <= 8'hbc;
      11'd1087 : out_data_ref <= 8'h6f;
      11'd1088 : out_data_ref <= 8'h96;
      11'd1089 : out_data_ref <= 8'h5b;
      11'd1090 : out_data_ref <= 8'h75;
      11'd1091 : out_data_ref <= 8'hfe;
      11'd1092 : out_data_ref <= 8'h59;
      11'd1093 : out_data_ref <= 8'ha5;
      11'd1094 : out_data_ref <= 8'haf;
      11'd1095 : out_data_ref <= 8'h29;
      11'd1096 : out_data_ref <= 8'h77;
      11'd1097 : out_data_ref <= 8'hd8;
      11'd1098 : out_data_ref <= 8'h1a;
      11'd1099 : out_data_ref <= 8'h0f;
      11'd1100 : out_data_ref <= 8'hb7;
      11'd1101 : out_data_ref <= 8'h33;
      11'd1102 : out_data_ref <= 8'h5d;
      11'd1103 : out_data_ref <= 8'h80;
      11'd1104 : out_data_ref <= 8'hac;
      11'd1105 : out_data_ref <= 8'h27;
      11'd1106 : out_data_ref <= 8'h68;
      11'd1107 : out_data_ref <= 8'hbf;
      11'd1108 : out_data_ref <= 8'h02;
      11'd1109 : out_data_ref <= 8'h2e;
      11'd1110 : out_data_ref <= 8'h27;
      11'd1111 : out_data_ref <= 8'hda;
      11'd1112 : out_data_ref <= 8'hc6;
      11'd1113 : out_data_ref <= 8'h6d;
      11'd1114 : out_data_ref <= 8'h21;
      11'd1115 : out_data_ref <= 8'h37;
      11'd1116 : out_data_ref <= 8'ha0;
      11'd1117 : out_data_ref <= 8'hb3;
      11'd1118 : out_data_ref <= 8'ha0;
      11'd1119 : out_data_ref <= 8'h7e;
      11'd1120 : out_data_ref <= 8'hdf;
      11'd1121 : out_data_ref <= 8'h71;
      11'd1122 : out_data_ref <= 8'h02;
      11'd1123 : out_data_ref <= 8'h21;
      11'd1124 : out_data_ref <= 8'h9d;
      11'd1125 : out_data_ref <= 8'h8c;
      11'd1126 : out_data_ref <= 8'h61;
      11'd1127 : out_data_ref <= 8'h98;
      11'd1128 : out_data_ref <= 8'hf0;
      11'd1129 : out_data_ref <= 8'h26;
      11'd1130 : out_data_ref <= 8'h3e;
      11'd1131 : out_data_ref <= 8'h35;
      11'd1132 : out_data_ref <= 8'h09;
      11'd1133 : out_data_ref <= 8'h3d;
      11'd1134 : out_data_ref <= 8'hfe;
      11'd1135 : out_data_ref <= 8'h97;
      11'd1136 : out_data_ref <= 8'hc2;
      11'd1137 : out_data_ref <= 8'hd8;
      11'd1138 : out_data_ref <= 8'hbb;
      11'd1139 : out_data_ref <= 8'h95;
      11'd1140 : out_data_ref <= 8'h79;
      11'd1141 : out_data_ref <= 8'h3f;
      11'd1142 : out_data_ref <= 8'hb9;
      11'd1143 : out_data_ref <= 8'h60;
      11'd1144 : out_data_ref <= 8'h23;
      11'd1145 : out_data_ref <= 8'hb6;
      11'd1146 : out_data_ref <= 8'he6;
      11'd1147 : out_data_ref <= 8'hdd;
      11'd1148 : out_data_ref <= 8'ha8;
      11'd1149 : out_data_ref <= 8'h5a;
      11'd1150 : out_data_ref <= 8'haa;
      11'd1151 : out_data_ref <= 8'hcf;
      11'd1152 : out_data_ref <= 8'h8b;
      11'd1153 : out_data_ref <= 8'h87;
      11'd1154 : out_data_ref <= 8'h39;
      11'd1155 : out_data_ref <= 8'h1b;
      11'd1156 : out_data_ref <= 8'h57;
      11'd1157 : out_data_ref <= 8'he9;
      11'd1158 : out_data_ref <= 8'hbc;
      11'd1159 : out_data_ref <= 8'h8c;
      11'd1160 : out_data_ref <= 8'hfe;
      11'd1161 : out_data_ref <= 8'h7f;
      11'd1162 : out_data_ref <= 8'he2;
      11'd1163 : out_data_ref <= 8'hd4;
      11'd1164 : out_data_ref <= 8'had;
      11'd1165 : out_data_ref <= 8'h98;
      11'd1166 : out_data_ref <= 8'h48;
      11'd1167 : out_data_ref <= 8'h7a;
      11'd1168 : out_data_ref <= 8'h79;
      11'd1169 : out_data_ref <= 8'h63;
      11'd1170 : out_data_ref <= 8'hcd;
      11'd1171 : out_data_ref <= 8'h9c;
      11'd1172 : out_data_ref <= 8'h0a;
      11'd1173 : out_data_ref <= 8'hd8;
      11'd1174 : out_data_ref <= 8'h0e;
      11'd1175 : out_data_ref <= 8'heb;
      11'd1176 : out_data_ref <= 8'h3b;
      11'd1177 : out_data_ref <= 8'h8c;
      11'd1178 : out_data_ref <= 8'h73;
      11'd1179 : out_data_ref <= 8'h12;
      11'd1180 : out_data_ref <= 8'h0d;
      11'd1181 : out_data_ref <= 8'hef;
      11'd1182 : out_data_ref <= 8'h03;
      11'd1183 : out_data_ref <= 8'hef;
      11'd1184 : out_data_ref <= 8'h3d;
      11'd1185 : out_data_ref <= 8'h3a;
      11'd1186 : out_data_ref <= 8'h43;
      11'd1187 : out_data_ref <= 8'hb1;
      11'd1188 : out_data_ref <= 8'h5d;
      11'd1189 : out_data_ref <= 8'h88;
      11'd1190 : out_data_ref <= 8'h08;
      11'd1191 : out_data_ref <= 8'hf8;
      11'd1192 : out_data_ref <= 8'ha7;
      11'd1193 : out_data_ref <= 8'h8d;
      11'd1194 : out_data_ref <= 8'h6a;
      11'd1195 : out_data_ref <= 8'h86;
      11'd1196 : out_data_ref <= 8'h7a;
      11'd1197 : out_data_ref <= 8'hd9;
      11'd1198 : out_data_ref <= 8'ha0;
      11'd1199 : out_data_ref <= 8'he8;
      11'd1200 : out_data_ref <= 8'h74;
      11'd1201 : out_data_ref <= 8'h47;
      11'd1202 : out_data_ref <= 8'hb8;
      11'd1203 : out_data_ref <= 8'hd2;
      11'd1204 : out_data_ref <= 8'h1b;
      11'd1205 : out_data_ref <= 8'he0;
      11'd1206 : out_data_ref <= 8'hc2;
      11'd1207 : out_data_ref <= 8'h7f;
      11'd1208 : out_data_ref <= 8'h30;
      11'd1209 : out_data_ref <= 8'ha1;
      11'd1210 : out_data_ref <= 8'hf5;
      11'd1211 : out_data_ref <= 8'ha2;
      11'd1212 : out_data_ref <= 8'h22;
      11'd1213 : out_data_ref <= 8'ha4;
      11'd1214 : out_data_ref <= 8'hac;
      11'd1215 : out_data_ref <= 8'h40;
      11'd1216 : out_data_ref <= 8'h2e;
      11'd1217 : out_data_ref <= 8'h57;
      11'd1218 : out_data_ref <= 8'h6c;
      11'd1219 : out_data_ref <= 8'hb9;
      11'd1220 : out_data_ref <= 8'h07;
      11'd1221 : out_data_ref <= 8'h84;
      11'd1222 : out_data_ref <= 8'hca;
      11'd1223 : out_data_ref <= 8'h05;
      11'd1224 : out_data_ref <= 8'hde;
      11'd1225 : out_data_ref <= 8'h12;
      11'd1226 : out_data_ref <= 8'hfd;
      11'd1227 : out_data_ref <= 8'hcf;
      11'd1228 : out_data_ref <= 8'he3;
      11'd1229 : out_data_ref <= 8'hee;
      11'd1230 : out_data_ref <= 8'h1e;
      11'd1231 : out_data_ref <= 8'h40;
      11'd1232 : out_data_ref <= 8'h71;
      11'd1233 : out_data_ref <= 8'hb9;
      11'd1234 : out_data_ref <= 8'h9d;
      11'd1235 : out_data_ref <= 8'h27;
      11'd1236 : out_data_ref <= 8'hf5;
      11'd1237 : out_data_ref <= 8'h14;
      11'd1238 : out_data_ref <= 8'h3c;
      11'd1239 : out_data_ref <= 8'h97;
      11'd1240 : out_data_ref <= 8'hd3;
      11'd1241 : out_data_ref <= 8'h03;
      11'd1242 : out_data_ref <= 8'ha5;
      11'd1243 : out_data_ref <= 8'h6a;
      11'd1244 : out_data_ref <= 8'h38;
      11'd1245 : out_data_ref <= 8'h7b;
      11'd1246 : out_data_ref <= 8'hfc;
      11'd1247 : out_data_ref <= 8'h4c;
      11'd1248 : out_data_ref <= 8'hb8;
      11'd1249 : out_data_ref <= 8'hcb;
      11'd1250 : out_data_ref <= 8'hdb;
      11'd1251 : out_data_ref <= 8'hbe;
      11'd1252 : out_data_ref <= 8'h0b;
      11'd1253 : out_data_ref <= 8'h68;
      11'd1254 : out_data_ref <= 8'hc4;
      11'd1255 : out_data_ref <= 8'h67;
      11'd1256 : out_data_ref <= 8'hca;
      11'd1257 : out_data_ref <= 8'h2c;
      11'd1258 : out_data_ref <= 8'h76;
      11'd1259 : out_data_ref <= 8'hdb;
      11'd1260 : out_data_ref <= 8'h00;
      11'd1261 : out_data_ref <= 8'h92;
      11'd1262 : out_data_ref <= 8'h6d;
      11'd1263 : out_data_ref <= 8'he2;
      11'd1264 : out_data_ref <= 8'h1d;
      11'd1265 : out_data_ref <= 8'h1f;
      11'd1266 : out_data_ref <= 8'h7d;
      11'd1267 : out_data_ref <= 8'h29;
      11'd1268 : out_data_ref <= 8'h09;
      11'd1269 : out_data_ref <= 8'h3e;
      11'd1270 : out_data_ref <= 8'h2f;
      11'd1271 : out_data_ref <= 8'hdc;
      11'd1272 : out_data_ref <= 8'hdd;
      11'd1273 : out_data_ref <= 8'ha9;
      11'd1274 : out_data_ref <= 8'h9c;
      11'd1275 : out_data_ref <= 8'hfb;
      11'd1276 : out_data_ref <= 8'h37;
      11'd1277 : out_data_ref <= 8'hd6;
      11'd1278 : out_data_ref <= 8'hb9;
      11'd1279 : out_data_ref <= 8'h9d;
      11'd1280 : out_data_ref <= 8'h6a;
      11'd1281 : out_data_ref <= 8'haf;
      11'd1282 : out_data_ref <= 8'hb3;
      11'd1283 : out_data_ref <= 8'h7d;
      11'd1284 : out_data_ref <= 8'hcd;
      11'd1285 : out_data_ref <= 8'hc6;
      11'd1286 : out_data_ref <= 8'h1f;
      11'd1287 : out_data_ref <= 8'h1f;
      11'd1288 : out_data_ref <= 8'h14;
      11'd1289 : out_data_ref <= 8'hba;
      11'd1290 : out_data_ref <= 8'h57;
      11'd1291 : out_data_ref <= 8'he3;
      11'd1292 : out_data_ref <= 8'h31;
      11'd1293 : out_data_ref <= 8'h76;
      11'd1294 : out_data_ref <= 8'h7d;
      11'd1295 : out_data_ref <= 8'h75;
      11'd1296 : out_data_ref <= 8'h07;
      11'd1297 : out_data_ref <= 8'he1;
      11'd1298 : out_data_ref <= 8'hc1;
      11'd1299 : out_data_ref <= 8'hc5;
      11'd1300 : out_data_ref <= 8'hdc;
      11'd1301 : out_data_ref <= 8'h54;
      11'd1302 : out_data_ref <= 8'h23;
      11'd1303 : out_data_ref <= 8'h49;
      11'd1304 : out_data_ref <= 8'hba;
      11'd1305 : out_data_ref <= 8'h23;
      11'd1306 : out_data_ref <= 8'h83;
      11'd1307 : out_data_ref <= 8'h6c;
      11'd1308 : out_data_ref <= 8'h71;
      11'd1309 : out_data_ref <= 8'hf4;
      11'd1310 : out_data_ref <= 8'he0;
      11'd1311 : out_data_ref <= 8'hfe;
      11'd1312 : out_data_ref <= 8'hc6;
      11'd1313 : out_data_ref <= 8'ha8;
      11'd1314 : out_data_ref <= 8'h13;
      11'd1315 : out_data_ref <= 8'hde;
      11'd1316 : out_data_ref <= 8'hd5;
      11'd1317 : out_data_ref <= 8'h9d;
      11'd1318 : out_data_ref <= 8'h14;
      11'd1319 : out_data_ref <= 8'ha2;
      11'd1320 : out_data_ref <= 8'h30;
      11'd1321 : out_data_ref <= 8'h10;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
