module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam B_LEN = 'd994;
  localparam B_DEPTH = 'd10;
  localparam R_LEN = 'd653;
  localparam R_DEPTH = 'd10;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [ 7: 0] in_data;
  input      [ 9: 0] out_addr;
  output reg [13: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 8'h01;
      10'd1    : in_data <= 8'h03;
      10'd2    : in_data <= 8'h1f;
      10'd3    : in_data <= 8'he0;
      10'd4    : in_data <= 8'hc4;
      10'd5    : in_data <= 8'h32;
      10'd6    : in_data <= 8'h8b;
      10'd7    : in_data <= 8'h95;
      10'd8    : in_data <= 8'h6e;
      10'd9    : in_data <= 8'h9a;
      10'd10   : in_data <= 8'hfa;
      10'd11   : in_data <= 8'h7b;
      10'd12   : in_data <= 8'h5d;
      10'd13   : in_data <= 8'h86;
      10'd14   : in_data <= 8'hde;
      10'd15   : in_data <= 8'h2c;
      10'd16   : in_data <= 8'hbf;
      10'd17   : in_data <= 8'h1f;
      10'd18   : in_data <= 8'h07;
      10'd19   : in_data <= 8'h28;
      10'd20   : in_data <= 8'ha1;
      10'd21   : in_data <= 8'h23;
      10'd22   : in_data <= 8'h6f;
      10'd23   : in_data <= 8'h68;
      10'd24   : in_data <= 8'h5d;
      10'd25   : in_data <= 8'hd2;
      10'd26   : in_data <= 8'hfd;
      10'd27   : in_data <= 8'h22;
      10'd28   : in_data <= 8'h1a;
      10'd29   : in_data <= 8'hcd;
      10'd30   : in_data <= 8'hd0;
      10'd31   : in_data <= 8'h5c;
      10'd32   : in_data <= 8'hab;
      10'd33   : in_data <= 8'h64;
      10'd34   : in_data <= 8'hb0;
      10'd35   : in_data <= 8'h1a;
      10'd36   : in_data <= 8'hf7;
      10'd37   : in_data <= 8'ha5;
      10'd38   : in_data <= 8'hf3;
      10'd39   : in_data <= 8'hc2;
      10'd40   : in_data <= 8'h83;
      10'd41   : in_data <= 8'h7a;
      10'd42   : in_data <= 8'h5b;
      10'd43   : in_data <= 8'h7f;
      10'd44   : in_data <= 8'he5;
      10'd45   : in_data <= 8'hfe;
      10'd46   : in_data <= 8'h31;
      10'd47   : in_data <= 8'he3;
      10'd48   : in_data <= 8'h66;
      10'd49   : in_data <= 8'hf7;
      10'd50   : in_data <= 8'hf0;
      10'd51   : in_data <= 8'h4c;
      10'd52   : in_data <= 8'h5b;
      10'd53   : in_data <= 8'h77;
      10'd54   : in_data <= 8'hc1;
      10'd55   : in_data <= 8'hd6;
      10'd56   : in_data <= 8'hbd;
      10'd57   : in_data <= 8'h3b;
      10'd58   : in_data <= 8'h25;
      10'd59   : in_data <= 8'ha7;
      10'd60   : in_data <= 8'h65;
      10'd61   : in_data <= 8'ha8;
      10'd62   : in_data <= 8'h4c;
      10'd63   : in_data <= 8'hf9;
      10'd64   : in_data <= 8'haa;
      10'd65   : in_data <= 8'h08;
      10'd66   : in_data <= 8'hfd;
      10'd67   : in_data <= 8'h9a;
      10'd68   : in_data <= 8'hba;
      10'd69   : in_data <= 8'h3b;
      10'd70   : in_data <= 8'hb6;
      10'd71   : in_data <= 8'ha4;
      10'd72   : in_data <= 8'hb5;
      10'd73   : in_data <= 8'hc3;
      10'd74   : in_data <= 8'h50;
      10'd75   : in_data <= 8'h40;
      10'd76   : in_data <= 8'h64;
      10'd77   : in_data <= 8'hd0;
      10'd78   : in_data <= 8'h80;
      10'd79   : in_data <= 8'h36;
      10'd80   : in_data <= 8'h87;
      10'd81   : in_data <= 8'ha0;
      10'd82   : in_data <= 8'h4f;
      10'd83   : in_data <= 8'h06;
      10'd84   : in_data <= 8'hb2;
      10'd85   : in_data <= 8'hbb;
      10'd86   : in_data <= 8'h5f;
      10'd87   : in_data <= 8'h7b;
      10'd88   : in_data <= 8'hb9;
      10'd89   : in_data <= 8'h5a;
      10'd90   : in_data <= 8'hab;
      10'd91   : in_data <= 8'hf6;
      10'd92   : in_data <= 8'hcb;
      10'd93   : in_data <= 8'h82;
      10'd94   : in_data <= 8'h3a;
      10'd95   : in_data <= 8'hcc;
      10'd96   : in_data <= 8'h6e;
      10'd97   : in_data <= 8'h74;
      10'd98   : in_data <= 8'he9;
      10'd99   : in_data <= 8'h8f;
      10'd100  : in_data <= 8'hc4;
      10'd101  : in_data <= 8'h68;
      10'd102  : in_data <= 8'hc3;
      10'd103  : in_data <= 8'he0;
      10'd104  : in_data <= 8'h7b;
      10'd105  : in_data <= 8'hca;
      10'd106  : in_data <= 8'he2;
      10'd107  : in_data <= 8'h84;
      10'd108  : in_data <= 8'h79;
      10'd109  : in_data <= 8'h72;
      10'd110  : in_data <= 8'h21;
      10'd111  : in_data <= 8'ha8;
      10'd112  : in_data <= 8'hc8;
      10'd113  : in_data <= 8'ha1;
      10'd114  : in_data <= 8'h61;
      10'd115  : in_data <= 8'h68;
      10'd116  : in_data <= 8'ha9;
      10'd117  : in_data <= 8'h1a;
      10'd118  : in_data <= 8'h03;
      10'd119  : in_data <= 8'hd0;
      10'd120  : in_data <= 8'h66;
      10'd121  : in_data <= 8'hf0;
      10'd122  : in_data <= 8'hec;
      10'd123  : in_data <= 8'h93;
      10'd124  : in_data <= 8'hf2;
      10'd125  : in_data <= 8'h6c;
      10'd126  : in_data <= 8'h8b;
      10'd127  : in_data <= 8'hb6;
      10'd128  : in_data <= 8'he9;
      10'd129  : in_data <= 8'h48;
      10'd130  : in_data <= 8'hbe;
      10'd131  : in_data <= 8'hcb;
      10'd132  : in_data <= 8'h99;
      10'd133  : in_data <= 8'h19;
      10'd134  : in_data <= 8'ha7;
      10'd135  : in_data <= 8'h2e;
      10'd136  : in_data <= 8'h0f;
      10'd137  : in_data <= 8'hb8;
      10'd138  : in_data <= 8'h6f;
      10'd139  : in_data <= 8'h38;
      10'd140  : in_data <= 8'h0f;
      10'd141  : in_data <= 8'h1f;
      10'd142  : in_data <= 8'h2c;
      10'd143  : in_data <= 8'h1a;
      10'd144  : in_data <= 8'h2e;
      10'd145  : in_data <= 8'hfc;
      10'd146  : in_data <= 8'hef;
      10'd147  : in_data <= 8'h87;
      10'd148  : in_data <= 8'h1d;
      10'd149  : in_data <= 8'h6a;
      10'd150  : in_data <= 8'hce;
      10'd151  : in_data <= 8'h4f;
      10'd152  : in_data <= 8'h5e;
      10'd153  : in_data <= 8'h0a;
      10'd154  : in_data <= 8'hd2;
      10'd155  : in_data <= 8'h26;
      10'd156  : in_data <= 8'ha8;
      10'd157  : in_data <= 8'h01;
      10'd158  : in_data <= 8'h17;
      10'd159  : in_data <= 8'hf7;
      10'd160  : in_data <= 8'hce;
      10'd161  : in_data <= 8'hef;
      10'd162  : in_data <= 8'he5;
      10'd163  : in_data <= 8'h66;
      10'd164  : in_data <= 8'h19;
      10'd165  : in_data <= 8'h3d;
      10'd166  : in_data <= 8'h87;
      10'd167  : in_data <= 8'h2a;
      10'd168  : in_data <= 8'h9a;
      10'd169  : in_data <= 8'hba;
      10'd170  : in_data <= 8'hdb;
      10'd171  : in_data <= 8'h98;
      10'd172  : in_data <= 8'h73;
      10'd173  : in_data <= 8'hd3;
      10'd174  : in_data <= 8'he9;
      10'd175  : in_data <= 8'hab;
      10'd176  : in_data <= 8'hb0;
      10'd177  : in_data <= 8'h11;
      10'd178  : in_data <= 8'h9c;
      10'd179  : in_data <= 8'hf4;
      10'd180  : in_data <= 8'h13;
      10'd181  : in_data <= 8'h3d;
      10'd182  : in_data <= 8'h06;
      10'd183  : in_data <= 8'hf0;
      10'd184  : in_data <= 8'hda;
      10'd185  : in_data <= 8'h9f;
      10'd186  : in_data <= 8'h0e;
      10'd187  : in_data <= 8'hcb;
      10'd188  : in_data <= 8'h63;
      10'd189  : in_data <= 8'h19;
      10'd190  : in_data <= 8'hce;
      10'd191  : in_data <= 8'he7;
      10'd192  : in_data <= 8'h96;
      10'd193  : in_data <= 8'hf2;
      10'd194  : in_data <= 8'hff;
      10'd195  : in_data <= 8'h5b;
      10'd196  : in_data <= 8'h85;
      10'd197  : in_data <= 8'hb4;
      10'd198  : in_data <= 8'ha6;
      10'd199  : in_data <= 8'h75;
      10'd200  : in_data <= 8'h4a;
      10'd201  : in_data <= 8'hd4;
      10'd202  : in_data <= 8'hc9;
      10'd203  : in_data <= 8'h43;
      10'd204  : in_data <= 8'h46;
      10'd205  : in_data <= 8'he3;
      10'd206  : in_data <= 8'h25;
      10'd207  : in_data <= 8'hba;
      10'd208  : in_data <= 8'hff;
      10'd209  : in_data <= 8'h9c;
      10'd210  : in_data <= 8'hc9;
      10'd211  : in_data <= 8'h22;
      10'd212  : in_data <= 8'h56;
      10'd213  : in_data <= 8'h1c;
      10'd214  : in_data <= 8'hf0;
      10'd215  : in_data <= 8'h2b;
      10'd216  : in_data <= 8'h82;
      10'd217  : in_data <= 8'h7e;
      10'd218  : in_data <= 8'h2a;
      10'd219  : in_data <= 8'h48;
      10'd220  : in_data <= 8'h7e;
      10'd221  : in_data <= 8'hce;
      10'd222  : in_data <= 8'h6a;
      10'd223  : in_data <= 8'h4a;
      10'd224  : in_data <= 8'hd9;
      10'd225  : in_data <= 8'hab;
      10'd226  : in_data <= 8'hbd;
      10'd227  : in_data <= 8'he1;
      10'd228  : in_data <= 8'hd8;
      10'd229  : in_data <= 8'h1c;
      10'd230  : in_data <= 8'h21;
      10'd231  : in_data <= 8'h8c;
      10'd232  : in_data <= 8'hd5;
      10'd233  : in_data <= 8'hd5;
      10'd234  : in_data <= 8'h0a;
      10'd235  : in_data <= 8'h66;
      10'd236  : in_data <= 8'hb8;
      10'd237  : in_data <= 8'he3;
      10'd238  : in_data <= 8'heb;
      10'd239  : in_data <= 8'h98;
      10'd240  : in_data <= 8'h70;
      10'd241  : in_data <= 8'hc9;
      10'd242  : in_data <= 8'hf6;
      10'd243  : in_data <= 8'h84;
      10'd244  : in_data <= 8'h57;
      10'd245  : in_data <= 8'hbc;
      10'd246  : in_data <= 8'h81;
      10'd247  : in_data <= 8'h3a;
      10'd248  : in_data <= 8'h2d;
      10'd249  : in_data <= 8'h82;
      10'd250  : in_data <= 8'h7e;
      10'd251  : in_data <= 8'ha7;
      10'd252  : in_data <= 8'hc8;
      10'd253  : in_data <= 8'h79;
      10'd254  : in_data <= 8'h51;
      10'd255  : in_data <= 8'h43;
      10'd256  : in_data <= 8'h9d;
      10'd257  : in_data <= 8'hd3;
      10'd258  : in_data <= 8'h94;
      10'd259  : in_data <= 8'hda;
      10'd260  : in_data <= 8'h1e;
      10'd261  : in_data <= 8'hd0;
      10'd262  : in_data <= 8'h71;
      10'd263  : in_data <= 8'he8;
      10'd264  : in_data <= 8'haa;
      10'd265  : in_data <= 8'hee;
      10'd266  : in_data <= 8'h17;
      10'd267  : in_data <= 8'h5b;
      10'd268  : in_data <= 8'hdb;
      10'd269  : in_data <= 8'hfc;
      10'd270  : in_data <= 8'h5c;
      10'd271  : in_data <= 8'he2;
      10'd272  : in_data <= 8'hac;
      10'd273  : in_data <= 8'hde;
      10'd274  : in_data <= 8'h12;
      10'd275  : in_data <= 8'hf7;
      10'd276  : in_data <= 8'h8c;
      10'd277  : in_data <= 8'h9b;
      10'd278  : in_data <= 8'h82;
      10'd279  : in_data <= 8'hd9;
      10'd280  : in_data <= 8'h65;
      10'd281  : in_data <= 8'h3b;
      10'd282  : in_data <= 8'h97;
      10'd283  : in_data <= 8'h0f;
      10'd284  : in_data <= 8'h03;
      10'd285  : in_data <= 8'h5a;
      10'd286  : in_data <= 8'h13;
      10'd287  : in_data <= 8'h0a;
      10'd288  : in_data <= 8'h1d;
      10'd289  : in_data <= 8'hfb;
      10'd290  : in_data <= 8'he5;
      10'd291  : in_data <= 8'hb2;
      10'd292  : in_data <= 8'hd4;
      10'd293  : in_data <= 8'hc1;
      10'd294  : in_data <= 8'h86;
      10'd295  : in_data <= 8'hc9;
      10'd296  : in_data <= 8'h09;
      10'd297  : in_data <= 8'hb9;
      10'd298  : in_data <= 8'had;
      10'd299  : in_data <= 8'hf4;
      10'd300  : in_data <= 8'hfb;
      10'd301  : in_data <= 8'h82;
      10'd302  : in_data <= 8'h1b;
      10'd303  : in_data <= 8'h2f;
      10'd304  : in_data <= 8'ha2;
      10'd305  : in_data <= 8'h1e;
      10'd306  : in_data <= 8'hc0;
      10'd307  : in_data <= 8'h3d;
      10'd308  : in_data <= 8'h8d;
      10'd309  : in_data <= 8'h8e;
      10'd310  : in_data <= 8'h09;
      10'd311  : in_data <= 8'h5d;
      10'd312  : in_data <= 8'h68;
      10'd313  : in_data <= 8'hf4;
      10'd314  : in_data <= 8'hcc;
      10'd315  : in_data <= 8'h12;
      10'd316  : in_data <= 8'hce;
      10'd317  : in_data <= 8'hdb;
      10'd318  : in_data <= 8'he1;
      10'd319  : in_data <= 8'hde;
      10'd320  : in_data <= 8'h74;
      10'd321  : in_data <= 8'h28;
      10'd322  : in_data <= 8'ha2;
      10'd323  : in_data <= 8'h01;
      10'd324  : in_data <= 8'hb0;
      10'd325  : in_data <= 8'h4a;
      10'd326  : in_data <= 8'h95;
      10'd327  : in_data <= 8'h75;
      10'd328  : in_data <= 8'hbe;
      10'd329  : in_data <= 8'h75;
      10'd330  : in_data <= 8'h8d;
      10'd331  : in_data <= 8'h58;
      10'd332  : in_data <= 8'h34;
      10'd333  : in_data <= 8'h0e;
      10'd334  : in_data <= 8'h73;
      10'd335  : in_data <= 8'h60;
      10'd336  : in_data <= 8'h2c;
      10'd337  : in_data <= 8'h34;
      10'd338  : in_data <= 8'h67;
      10'd339  : in_data <= 8'h87;
      10'd340  : in_data <= 8'h6a;
      10'd341  : in_data <= 8'h4b;
      10'd342  : in_data <= 8'h18;
      10'd343  : in_data <= 8'h21;
      10'd344  : in_data <= 8'h8c;
      10'd345  : in_data <= 8'h34;
      10'd346  : in_data <= 8'ha3;
      10'd347  : in_data <= 8'h12;
      10'd348  : in_data <= 8'h6d;
      10'd349  : in_data <= 8'hbc;
      10'd350  : in_data <= 8'hc8;
      10'd351  : in_data <= 8'h77;
      10'd352  : in_data <= 8'h14;
      10'd353  : in_data <= 8'h4e;
      10'd354  : in_data <= 8'h4a;
      10'd355  : in_data <= 8'h42;
      10'd356  : in_data <= 8'ha4;
      10'd357  : in_data <= 8'h50;
      10'd358  : in_data <= 8'h05;
      10'd359  : in_data <= 8'h21;
      10'd360  : in_data <= 8'h7d;
      10'd361  : in_data <= 8'h9c;
      10'd362  : in_data <= 8'h50;
      10'd363  : in_data <= 8'hf3;
      10'd364  : in_data <= 8'h8d;
      10'd365  : in_data <= 8'hba;
      10'd366  : in_data <= 8'hfa;
      10'd367  : in_data <= 8'hc6;
      10'd368  : in_data <= 8'h47;
      10'd369  : in_data <= 8'h70;
      10'd370  : in_data <= 8'h11;
      10'd371  : in_data <= 8'hda;
      10'd372  : in_data <= 8'h1a;
      10'd373  : in_data <= 8'h1f;
      10'd374  : in_data <= 8'hc7;
      10'd375  : in_data <= 8'h49;
      10'd376  : in_data <= 8'hf2;
      10'd377  : in_data <= 8'h6b;
      10'd378  : in_data <= 8'h6c;
      10'd379  : in_data <= 8'h74;
      10'd380  : in_data <= 8'h7d;
      10'd381  : in_data <= 8'hda;
      10'd382  : in_data <= 8'hdf;
      10'd383  : in_data <= 8'h1f;
      10'd384  : in_data <= 8'h1e;
      10'd385  : in_data <= 8'h47;
      10'd386  : in_data <= 8'h07;
      10'd387  : in_data <= 8'h44;
      10'd388  : in_data <= 8'h0a;
      10'd389  : in_data <= 8'h34;
      10'd390  : in_data <= 8'hc2;
      10'd391  : in_data <= 8'h20;
      10'd392  : in_data <= 8'h46;
      10'd393  : in_data <= 8'ha6;
      10'd394  : in_data <= 8'h14;
      10'd395  : in_data <= 8'h5d;
      10'd396  : in_data <= 8'h30;
      10'd397  : in_data <= 8'h33;
      10'd398  : in_data <= 8'h40;
      10'd399  : in_data <= 8'h82;
      10'd400  : in_data <= 8'h12;
      10'd401  : in_data <= 8'h25;
      10'd402  : in_data <= 8'h4f;
      10'd403  : in_data <= 8'hbe;
      10'd404  : in_data <= 8'hfa;
      10'd405  : in_data <= 8'he6;
      10'd406  : in_data <= 8'ha4;
      10'd407  : in_data <= 8'hfc;
      10'd408  : in_data <= 8'hf5;
      10'd409  : in_data <= 8'haa;
      10'd410  : in_data <= 8'h41;
      10'd411  : in_data <= 8'hba;
      10'd412  : in_data <= 8'h14;
      10'd413  : in_data <= 8'hef;
      10'd414  : in_data <= 8'h3c;
      10'd415  : in_data <= 8'h6c;
      10'd416  : in_data <= 8'ha2;
      10'd417  : in_data <= 8'h3f;
      10'd418  : in_data <= 8'h3e;
      10'd419  : in_data <= 8'h04;
      10'd420  : in_data <= 8'hca;
      10'd421  : in_data <= 8'h53;
      10'd422  : in_data <= 8'ha5;
      10'd423  : in_data <= 8'hc2;
      10'd424  : in_data <= 8'haa;
      10'd425  : in_data <= 8'h03;
      10'd426  : in_data <= 8'hc7;
      10'd427  : in_data <= 8'h17;
      10'd428  : in_data <= 8'ha0;
      10'd429  : in_data <= 8'h4e;
      10'd430  : in_data <= 8'h92;
      10'd431  : in_data <= 8'h8e;
      10'd432  : in_data <= 8'h5d;
      10'd433  : in_data <= 8'hd3;
      10'd434  : in_data <= 8'h92;
      10'd435  : in_data <= 8'had;
      10'd436  : in_data <= 8'hfb;
      10'd437  : in_data <= 8'ha9;
      10'd438  : in_data <= 8'h21;
      10'd439  : in_data <= 8'h52;
      10'd440  : in_data <= 8'h8e;
      10'd441  : in_data <= 8'h54;
      10'd442  : in_data <= 8'h94;
      10'd443  : in_data <= 8'h4b;
      10'd444  : in_data <= 8'h41;
      10'd445  : in_data <= 8'h83;
      10'd446  : in_data <= 8'hac;
      10'd447  : in_data <= 8'hbe;
      10'd448  : in_data <= 8'hd4;
      10'd449  : in_data <= 8'hd2;
      10'd450  : in_data <= 8'h1d;
      10'd451  : in_data <= 8'hff;
      10'd452  : in_data <= 8'ha3;
      10'd453  : in_data <= 8'hf3;
      10'd454  : in_data <= 8'h3d;
      10'd455  : in_data <= 8'h35;
      10'd456  : in_data <= 8'hb9;
      10'd457  : in_data <= 8'h67;
      10'd458  : in_data <= 8'h90;
      10'd459  : in_data <= 8'h68;
      10'd460  : in_data <= 8'hb3;
      10'd461  : in_data <= 8'h71;
      10'd462  : in_data <= 8'h1a;
      10'd463  : in_data <= 8'hc4;
      10'd464  : in_data <= 8'h38;
      10'd465  : in_data <= 8'hf7;
      10'd466  : in_data <= 8'hca;
      10'd467  : in_data <= 8'hf3;
      10'd468  : in_data <= 8'h04;
      10'd469  : in_data <= 8'h24;
      10'd470  : in_data <= 8'h36;
      10'd471  : in_data <= 8'ha9;
      10'd472  : in_data <= 8'hc0;
      10'd473  : in_data <= 8'hbb;
      10'd474  : in_data <= 8'h29;
      10'd475  : in_data <= 8'h6e;
      10'd476  : in_data <= 8'hd1;
      10'd477  : in_data <= 8'hc7;
      10'd478  : in_data <= 8'h89;
      10'd479  : in_data <= 8'h1b;
      10'd480  : in_data <= 8'h7b;
      10'd481  : in_data <= 8'h78;
      10'd482  : in_data <= 8'h2e;
      10'd483  : in_data <= 8'haa;
      10'd484  : in_data <= 8'hbf;
      10'd485  : in_data <= 8'hce;
      10'd486  : in_data <= 8'h08;
      10'd487  : in_data <= 8'h0b;
      10'd488  : in_data <= 8'hdc;
      10'd489  : in_data <= 8'h54;
      10'd490  : in_data <= 8'hcb;
      10'd491  : in_data <= 8'h4e;
      10'd492  : in_data <= 8'hae;
      10'd493  : in_data <= 8'h3e;
      10'd494  : in_data <= 8'h75;
      10'd495  : in_data <= 8'h53;
      10'd496  : in_data <= 8'h61;
      10'd497  : in_data <= 8'h71;
      10'd498  : in_data <= 8'hbf;
      10'd499  : in_data <= 8'h12;
      10'd500  : in_data <= 8'h35;
      10'd501  : in_data <= 8'h39;
      10'd502  : in_data <= 8'h7e;
      10'd503  : in_data <= 8'hd3;
      10'd504  : in_data <= 8'h7a;
      10'd505  : in_data <= 8'h43;
      10'd506  : in_data <= 8'h94;
      10'd507  : in_data <= 8'hd0;
      10'd508  : in_data <= 8'h5d;
      10'd509  : in_data <= 8'h31;
      10'd510  : in_data <= 8'hd7;
      10'd511  : in_data <= 8'h27;
      10'd512  : in_data <= 8'h4a;
      10'd513  : in_data <= 8'h16;
      10'd514  : in_data <= 8'h40;
      10'd515  : in_data <= 8'hc1;
      10'd516  : in_data <= 8'hb4;
      10'd517  : in_data <= 8'h29;
      10'd518  : in_data <= 8'h12;
      10'd519  : in_data <= 8'hcd;
      10'd520  : in_data <= 8'h9a;
      10'd521  : in_data <= 8'heb;
      10'd522  : in_data <= 8'hb6;
      10'd523  : in_data <= 8'hb3;
      10'd524  : in_data <= 8'h23;
      10'd525  : in_data <= 8'hc3;
      10'd526  : in_data <= 8'h70;
      10'd527  : in_data <= 8'h13;
      10'd528  : in_data <= 8'h0a;
      10'd529  : in_data <= 8'h85;
      10'd530  : in_data <= 8'h4e;
      10'd531  : in_data <= 8'h5b;
      10'd532  : in_data <= 8'hb2;
      10'd533  : in_data <= 8'h25;
      10'd534  : in_data <= 8'h3d;
      10'd535  : in_data <= 8'h6f;
      10'd536  : in_data <= 8'h3c;
      10'd537  : in_data <= 8'ha7;
      10'd538  : in_data <= 8'haf;
      10'd539  : in_data <= 8'ha0;
      10'd540  : in_data <= 8'h61;
      10'd541  : in_data <= 8'hc2;
      10'd542  : in_data <= 8'h41;
      10'd543  : in_data <= 8'h64;
      10'd544  : in_data <= 8'h6c;
      10'd545  : in_data <= 8'h28;
      10'd546  : in_data <= 8'ha8;
      10'd547  : in_data <= 8'hd1;
      10'd548  : in_data <= 8'hea;
      10'd549  : in_data <= 8'h7a;
      10'd550  : in_data <= 8'hac;
      10'd551  : in_data <= 8'ha7;
      10'd552  : in_data <= 8'h3a;
      10'd553  : in_data <= 8'h02;
      10'd554  : in_data <= 8'h89;
      10'd555  : in_data <= 8'h20;
      10'd556  : in_data <= 8'hc2;
      10'd557  : in_data <= 8'hba;
      10'd558  : in_data <= 8'h5d;
      10'd559  : in_data <= 8'hc9;
      10'd560  : in_data <= 8'hec;
      10'd561  : in_data <= 8'h21;
      10'd562  : in_data <= 8'hf1;
      10'd563  : in_data <= 8'h64;
      10'd564  : in_data <= 8'h5b;
      10'd565  : in_data <= 8'h92;
      10'd566  : in_data <= 8'hb3;
      10'd567  : in_data <= 8'h5f;
      10'd568  : in_data <= 8'he8;
      10'd569  : in_data <= 8'h10;
      10'd570  : in_data <= 8'he0;
      10'd571  : in_data <= 8'h24;
      10'd572  : in_data <= 8'hcb;
      10'd573  : in_data <= 8'h76;
      10'd574  : in_data <= 8'h4c;
      10'd575  : in_data <= 8'he5;
      10'd576  : in_data <= 8'h3f;
      10'd577  : in_data <= 8'h61;
      10'd578  : in_data <= 8'h1e;
      10'd579  : in_data <= 8'h61;
      10'd580  : in_data <= 8'hdf;
      10'd581  : in_data <= 8'hc6;
      10'd582  : in_data <= 8'h2c;
      10'd583  : in_data <= 8'hed;
      10'd584  : in_data <= 8'hd8;
      10'd585  : in_data <= 8'hbc;
      10'd586  : in_data <= 8'hd4;
      10'd587  : in_data <= 8'h45;
      10'd588  : in_data <= 8'h87;
      10'd589  : in_data <= 8'h0d;
      10'd590  : in_data <= 8'h50;
      10'd591  : in_data <= 8'heb;
      10'd592  : in_data <= 8'hd4;
      10'd593  : in_data <= 8'hdd;
      10'd594  : in_data <= 8'h80;
      10'd595  : in_data <= 8'h21;
      10'd596  : in_data <= 8'h92;
      10'd597  : in_data <= 8'h4c;
      10'd598  : in_data <= 8'hc3;
      10'd599  : in_data <= 8'h66;
      10'd600  : in_data <= 8'hfa;
      10'd601  : in_data <= 8'hde;
      10'd602  : in_data <= 8'h33;
      10'd603  : in_data <= 8'h0a;
      10'd604  : in_data <= 8'hc3;
      10'd605  : in_data <= 8'h82;
      10'd606  : in_data <= 8'h6d;
      10'd607  : in_data <= 8'hbf;
      10'd608  : in_data <= 8'h43;
      10'd609  : in_data <= 8'ha3;
      10'd610  : in_data <= 8'h28;
      10'd611  : in_data <= 8'h25;
      10'd612  : in_data <= 8'h4c;
      10'd613  : in_data <= 8'h36;
      10'd614  : in_data <= 8'h7b;
      10'd615  : in_data <= 8'h15;
      10'd616  : in_data <= 8'h71;
      10'd617  : in_data <= 8'h89;
      10'd618  : in_data <= 8'h67;
      10'd619  : in_data <= 8'hd7;
      10'd620  : in_data <= 8'h2e;
      10'd621  : in_data <= 8'hb4;
      10'd622  : in_data <= 8'hf7;
      10'd623  : in_data <= 8'hec;
      10'd624  : in_data <= 8'h3b;
      10'd625  : in_data <= 8'hfb;
      10'd626  : in_data <= 8'h69;
      10'd627  : in_data <= 8'h2b;
      10'd628  : in_data <= 8'h5b;
      10'd629  : in_data <= 8'hef;
      10'd630  : in_data <= 8'h35;
      10'd631  : in_data <= 8'h7b;
      10'd632  : in_data <= 8'hef;
      10'd633  : in_data <= 8'h09;
      10'd634  : in_data <= 8'h74;
      10'd635  : in_data <= 8'h73;
      10'd636  : in_data <= 8'h94;
      10'd637  : in_data <= 8'h00;
      10'd638  : in_data <= 8'h11;
      10'd639  : in_data <= 8'h3f;
      10'd640  : in_data <= 8'h76;
      10'd641  : in_data <= 8'h69;
      10'd642  : in_data <= 8'h22;
      10'd643  : in_data <= 8'hf3;
      10'd644  : in_data <= 8'h17;
      10'd645  : in_data <= 8'h19;
      10'd646  : in_data <= 8'h64;
      10'd647  : in_data <= 8'he3;
      10'd648  : in_data <= 8'h03;
      10'd649  : in_data <= 8'hd2;
      10'd650  : in_data <= 8'h55;
      10'd651  : in_data <= 8'hfe;
      10'd652  : in_data <= 8'h24;
      10'd653  : in_data <= 8'h53;
      10'd654  : in_data <= 8'hbe;
      10'd655  : in_data <= 8'h85;
      10'd656  : in_data <= 8'haa;
      10'd657  : in_data <= 8'h7b;
      10'd658  : in_data <= 8'h9b;
      10'd659  : in_data <= 8'h9b;
      10'd660  : in_data <= 8'h64;
      10'd661  : in_data <= 8'h08;
      10'd662  : in_data <= 8'hd1;
      10'd663  : in_data <= 8'h65;
      10'd664  : in_data <= 8'h5d;
      10'd665  : in_data <= 8'h47;
      10'd666  : in_data <= 8'h5b;
      10'd667  : in_data <= 8'he7;
      10'd668  : in_data <= 8'hef;
      10'd669  : in_data <= 8'h03;
      10'd670  : in_data <= 8'h51;
      10'd671  : in_data <= 8'h27;
      10'd672  : in_data <= 8'h3b;
      10'd673  : in_data <= 8'hc0;
      10'd674  : in_data <= 8'h84;
      10'd675  : in_data <= 8'hc9;
      10'd676  : in_data <= 8'he7;
      10'd677  : in_data <= 8'h1b;
      10'd678  : in_data <= 8'h79;
      10'd679  : in_data <= 8'h4f;
      10'd680  : in_data <= 8'hac;
      10'd681  : in_data <= 8'h5c;
      10'd682  : in_data <= 8'h25;
      10'd683  : in_data <= 8'h6e;
      10'd684  : in_data <= 8'h87;
      10'd685  : in_data <= 8'hcf;
      10'd686  : in_data <= 8'hed;
      10'd687  : in_data <= 8'he5;
      10'd688  : in_data <= 8'hfd;
      10'd689  : in_data <= 8'h8e;
      10'd690  : in_data <= 8'h03;
      10'd691  : in_data <= 8'hec;
      10'd692  : in_data <= 8'h27;
      10'd693  : in_data <= 8'h2b;
      10'd694  : in_data <= 8'h24;
      10'd695  : in_data <= 8'h67;
      10'd696  : in_data <= 8'h5b;
      10'd697  : in_data <= 8'h94;
      10'd698  : in_data <= 8'h7b;
      10'd699  : in_data <= 8'hb5;
      10'd700  : in_data <= 8'hc1;
      10'd701  : in_data <= 8'h71;
      10'd702  : in_data <= 8'h1d;
      10'd703  : in_data <= 8'h89;
      10'd704  : in_data <= 8'h42;
      10'd705  : in_data <= 8'h85;
      10'd706  : in_data <= 8'he0;
      10'd707  : in_data <= 8'h26;
      10'd708  : in_data <= 8'h22;
      10'd709  : in_data <= 8'h1a;
      10'd710  : in_data <= 8'h15;
      10'd711  : in_data <= 8'h2d;
      10'd712  : in_data <= 8'h19;
      10'd713  : in_data <= 8'hdd;
      10'd714  : in_data <= 8'he6;
      10'd715  : in_data <= 8'h5e;
      10'd716  : in_data <= 8'hd2;
      10'd717  : in_data <= 8'h93;
      10'd718  : in_data <= 8'h71;
      10'd719  : in_data <= 8'h0d;
      10'd720  : in_data <= 8'h19;
      10'd721  : in_data <= 8'h5d;
      10'd722  : in_data <= 8'h31;
      10'd723  : in_data <= 8'h96;
      10'd724  : in_data <= 8'h8d;
      10'd725  : in_data <= 8'h18;
      10'd726  : in_data <= 8'he9;
      10'd727  : in_data <= 8'he2;
      10'd728  : in_data <= 8'hac;
      10'd729  : in_data <= 8'hf3;
      10'd730  : in_data <= 8'ha0;
      10'd731  : in_data <= 8'hbf;
      10'd732  : in_data <= 8'h5c;
      10'd733  : in_data <= 8'h9f;
      10'd734  : in_data <= 8'h47;
      10'd735  : in_data <= 8'h60;
      10'd736  : in_data <= 8'hb1;
      10'd737  : in_data <= 8'hc2;
      10'd738  : in_data <= 8'h0d;
      10'd739  : in_data <= 8'hdc;
      10'd740  : in_data <= 8'hb4;
      10'd741  : in_data <= 8'h9f;
      10'd742  : in_data <= 8'hd9;
      10'd743  : in_data <= 8'ha2;
      10'd744  : in_data <= 8'h4a;
      10'd745  : in_data <= 8'h30;
      10'd746  : in_data <= 8'h27;
      10'd747  : in_data <= 8'h02;
      10'd748  : in_data <= 8'h5a;
      10'd749  : in_data <= 8'h5c;
      10'd750  : in_data <= 8'h09;
      10'd751  : in_data <= 8'h0c;
      10'd752  : in_data <= 8'h70;
      10'd753  : in_data <= 8'h8e;
      10'd754  : in_data <= 8'h97;
      10'd755  : in_data <= 8'hcd;
      10'd756  : in_data <= 8'h0f;
      10'd757  : in_data <= 8'h27;
      10'd758  : in_data <= 8'h3e;
      10'd759  : in_data <= 8'h89;
      10'd760  : in_data <= 8'hdd;
      10'd761  : in_data <= 8'h43;
      10'd762  : in_data <= 8'h18;
      10'd763  : in_data <= 8'h0a;
      10'd764  : in_data <= 8'hbe;
      10'd765  : in_data <= 8'hac;
      10'd766  : in_data <= 8'h46;
      10'd767  : in_data <= 8'h65;
      10'd768  : in_data <= 8'h47;
      10'd769  : in_data <= 8'h87;
      10'd770  : in_data <= 8'h32;
      10'd771  : in_data <= 8'h68;
      10'd772  : in_data <= 8'h33;
      10'd773  : in_data <= 8'h25;
      10'd774  : in_data <= 8'h40;
      10'd775  : in_data <= 8'h6c;
      10'd776  : in_data <= 8'hfb;
      10'd777  : in_data <= 8'hf2;
      10'd778  : in_data <= 8'h0b;
      10'd779  : in_data <= 8'hf3;
      10'd780  : in_data <= 8'h05;
      10'd781  : in_data <= 8'h9a;
      10'd782  : in_data <= 8'he5;
      10'd783  : in_data <= 8'h77;
      10'd784  : in_data <= 8'h56;
      10'd785  : in_data <= 8'hfa;
      10'd786  : in_data <= 8'hf1;
      10'd787  : in_data <= 8'h85;
      10'd788  : in_data <= 8'h61;
      10'd789  : in_data <= 8'h2e;
      10'd790  : in_data <= 8'hc1;
      10'd791  : in_data <= 8'h99;
      10'd792  : in_data <= 8'h42;
      10'd793  : in_data <= 8'h4e;
      10'd794  : in_data <= 8'hc6;
      10'd795  : in_data <= 8'h4e;
      10'd796  : in_data <= 8'hc4;
      10'd797  : in_data <= 8'h44;
      10'd798  : in_data <= 8'hbc;
      10'd799  : in_data <= 8'h19;
      10'd800  : in_data <= 8'h0f;
      10'd801  : in_data <= 8'h0f;
      10'd802  : in_data <= 8'haa;
      10'd803  : in_data <= 8'h6b;
      10'd804  : in_data <= 8'h2e;
      10'd805  : in_data <= 8'h9a;
      10'd806  : in_data <= 8'h2d;
      10'd807  : in_data <= 8'h96;
      10'd808  : in_data <= 8'he7;
      10'd809  : in_data <= 8'h81;
      10'd810  : in_data <= 8'h4e;
      10'd811  : in_data <= 8'h2f;
      10'd812  : in_data <= 8'hc3;
      10'd813  : in_data <= 8'hbf;
      10'd814  : in_data <= 8'h67;
      10'd815  : in_data <= 8'h3b;
      10'd816  : in_data <= 8'h87;
      10'd817  : in_data <= 8'hb7;
      10'd818  : in_data <= 8'hce;
      10'd819  : in_data <= 8'hc8;
      10'd820  : in_data <= 8'hd6;
      10'd821  : in_data <= 8'hf3;
      10'd822  : in_data <= 8'ha8;
      10'd823  : in_data <= 8'h14;
      10'd824  : in_data <= 8'hb5;
      10'd825  : in_data <= 8'h77;
      10'd826  : in_data <= 8'h4c;
      10'd827  : in_data <= 8'hf9;
      10'd828  : in_data <= 8'h54;
      10'd829  : in_data <= 8'h90;
      10'd830  : in_data <= 8'he2;
      10'd831  : in_data <= 8'h58;
      10'd832  : in_data <= 8'hf0;
      10'd833  : in_data <= 8'hb1;
      10'd834  : in_data <= 8'h02;
      10'd835  : in_data <= 8'h69;
      10'd836  : in_data <= 8'he1;
      10'd837  : in_data <= 8'had;
      10'd838  : in_data <= 8'hd8;
      10'd839  : in_data <= 8'hc1;
      10'd840  : in_data <= 8'hd1;
      10'd841  : in_data <= 8'hc4;
      10'd842  : in_data <= 8'hbd;
      10'd843  : in_data <= 8'hd5;
      10'd844  : in_data <= 8'h34;
      10'd845  : in_data <= 8'h6a;
      10'd846  : in_data <= 8'hbd;
      10'd847  : in_data <= 8'h92;
      10'd848  : in_data <= 8'h1c;
      10'd849  : in_data <= 8'he3;
      10'd850  : in_data <= 8'he0;
      10'd851  : in_data <= 8'h2a;
      10'd852  : in_data <= 8'h2d;
      10'd853  : in_data <= 8'h05;
      10'd854  : in_data <= 8'h1a;
      10'd855  : in_data <= 8'h95;
      10'd856  : in_data <= 8'he5;
      10'd857  : in_data <= 8'h6d;
      10'd858  : in_data <= 8'hfe;
      10'd859  : in_data <= 8'h9a;
      10'd860  : in_data <= 8'h0c;
      10'd861  : in_data <= 8'h65;
      10'd862  : in_data <= 8'h5d;
      10'd863  : in_data <= 8'h92;
      10'd864  : in_data <= 8'h6f;
      10'd865  : in_data <= 8'hca;
      10'd866  : in_data <= 8'h45;
      10'd867  : in_data <= 8'hd4;
      10'd868  : in_data <= 8'h45;
      10'd869  : in_data <= 8'h17;
      10'd870  : in_data <= 8'h04;
      10'd871  : in_data <= 8'h98;
      10'd872  : in_data <= 8'hf6;
      10'd873  : in_data <= 8'hd0;
      10'd874  : in_data <= 8'h87;
      10'd875  : in_data <= 8'h0b;
      10'd876  : in_data <= 8'hc8;
      10'd877  : in_data <= 8'hd3;
      10'd878  : in_data <= 8'hf4;
      10'd879  : in_data <= 8'h44;
      10'd880  : in_data <= 8'h98;
      10'd881  : in_data <= 8'h2e;
      10'd882  : in_data <= 8'h55;
      10'd883  : in_data <= 8'hde;
      10'd884  : in_data <= 8'h23;
      10'd885  : in_data <= 8'hd5;
      10'd886  : in_data <= 8'h9a;
      10'd887  : in_data <= 8'h38;
      10'd888  : in_data <= 8'h5e;
      10'd889  : in_data <= 8'h1f;
      10'd890  : in_data <= 8'h18;
      10'd891  : in_data <= 8'h73;
      10'd892  : in_data <= 8'h2f;
      10'd893  : in_data <= 8'h7d;
      10'd894  : in_data <= 8'h7f;
      10'd895  : in_data <= 8'h65;
      10'd896  : in_data <= 8'h26;
      10'd897  : in_data <= 8'h28;
      10'd898  : in_data <= 8'h9c;
      10'd899  : in_data <= 8'h66;
      10'd900  : in_data <= 8'h59;
      10'd901  : in_data <= 8'hd4;
      10'd902  : in_data <= 8'h36;
      10'd903  : in_data <= 8'h30;
      10'd904  : in_data <= 8'h09;
      10'd905  : in_data <= 8'heb;
      10'd906  : in_data <= 8'hcd;
      10'd907  : in_data <= 8'hf2;
      10'd908  : in_data <= 8'h06;
      10'd909  : in_data <= 8'h64;
      10'd910  : in_data <= 8'h11;
      10'd911  : in_data <= 8'he4;
      10'd912  : in_data <= 8'h9e;
      10'd913  : in_data <= 8'h3a;
      10'd914  : in_data <= 8'h8e;
      10'd915  : in_data <= 8'h3d;
      10'd916  : in_data <= 8'h6b;
      10'd917  : in_data <= 8'h31;
      10'd918  : in_data <= 8'h2d;
      10'd919  : in_data <= 8'hdc;
      10'd920  : in_data <= 8'hc4;
      10'd921  : in_data <= 8'h91;
      10'd922  : in_data <= 8'h69;
      10'd923  : in_data <= 8'hbb;
      10'd924  : in_data <= 8'hf9;
      10'd925  : in_data <= 8'hb1;
      10'd926  : in_data <= 8'h3c;
      10'd927  : in_data <= 8'h82;
      10'd928  : in_data <= 8'h7a;
      10'd929  : in_data <= 8'h88;
      10'd930  : in_data <= 8'hac;
      10'd931  : in_data <= 8'hfd;
      10'd932  : in_data <= 8'h5b;
      10'd933  : in_data <= 8'h3e;
      10'd934  : in_data <= 8'h61;
      10'd935  : in_data <= 8'ha9;
      10'd936  : in_data <= 8'h11;
      10'd937  : in_data <= 8'h69;
      10'd938  : in_data <= 8'h16;
      10'd939  : in_data <= 8'hf4;
      10'd940  : in_data <= 8'h10;
      10'd941  : in_data <= 8'h52;
      10'd942  : in_data <= 8'ha3;
      10'd943  : in_data <= 8'haa;
      10'd944  : in_data <= 8'hf5;
      10'd945  : in_data <= 8'h0a;
      10'd946  : in_data <= 8'hbd;
      10'd947  : in_data <= 8'ha2;
      10'd948  : in_data <= 8'he7;
      10'd949  : in_data <= 8'hca;
      10'd950  : in_data <= 8'ha9;
      10'd951  : in_data <= 8'hdb;
      10'd952  : in_data <= 8'h7e;
      10'd953  : in_data <= 8'ha8;
      10'd954  : in_data <= 8'h16;
      10'd955  : in_data <= 8'hf4;
      10'd956  : in_data <= 8'h4c;
      10'd957  : in_data <= 8'h0f;
      10'd958  : in_data <= 8'h31;
      10'd959  : in_data <= 8'h5c;
      10'd960  : in_data <= 8'hb8;
      10'd961  : in_data <= 8'h67;
      10'd962  : in_data <= 8'h00;
      10'd963  : in_data <= 8'hf6;
      10'd964  : in_data <= 8'h2e;
      10'd965  : in_data <= 8'h25;
      10'd966  : in_data <= 8'he0;
      10'd967  : in_data <= 8'h5c;
      10'd968  : in_data <= 8'h90;
      10'd969  : in_data <= 8'h29;
      10'd970  : in_data <= 8'h4f;
      10'd971  : in_data <= 8'hbd;
      10'd972  : in_data <= 8'h55;
      10'd973  : in_data <= 8'h34;
      10'd974  : in_data <= 8'h2d;
      10'd975  : in_data <= 8'h62;
      10'd976  : in_data <= 8'hba;
      10'd977  : in_data <= 8'hfa;
      10'd978  : in_data <= 8'h8b;
      10'd979  : in_data <= 8'ha5;
      10'd980  : in_data <= 8'h5b;
      10'd981  : in_data <= 8'hee;
      10'd982  : in_data <= 8'h7b;
      10'd983  : in_data <= 8'h53;
      10'd984  : in_data <= 8'h2d;
      10'd985  : in_data <= 8'h50;
      10'd986  : in_data <= 8'hcd;
      10'd987  : in_data <= 8'h94;
      10'd988  : in_data <= 8'h70;
      10'd989  : in_data <= 8'h65;
      10'd990  : in_data <= 8'he7;
      10'd991  : in_data <= 8'h04;
      10'd992  : in_data <= 8'he6;
      10'd993  : in_data <= 8'h25;
      default: in_data <= 8'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      10'd0    : out_data_ref <= 14'h0a5d; // 'd2653
      10'd1    : out_data_ref <= 14'h0634; // 'd1588
      10'd2    : out_data_ref <= 14'h0fa7; // 'd4007
      10'd3    : out_data_ref <= 14'h0c58; // 'd3160
      10'd4    : out_data_ref <= 14'h076b; // 'd1899
      10'd5    : out_data_ref <= 14'h077d; // 'd1917
      10'd6    : out_data_ref <= 14'h028d; // 'd653
      10'd7    : out_data_ref <= 14'h0576; // 'd1398
      10'd8    : out_data_ref <= 14'h0549; // 'd1353
      10'd9    : out_data_ref <= 14'h0179; // 'd377
      10'd10   : out_data_ref <= 14'h115b; // 'd4443
      10'd11   : out_data_ref <= 14'h005b; // 'd91
      10'd12   : out_data_ref <= 14'h11e9; // 'd4585
      10'd13   : out_data_ref <= 14'h0d44; // 'd3396
      10'd14   : out_data_ref <= 14'h0384; // 'd900
      10'd15   : out_data_ref <= 14'h0a42; // 'd2626
      10'd16   : out_data_ref <= 14'h0460; // 'd1120
      10'd17   : out_data_ref <= 14'h041b; // 'd1051
      10'd18   : out_data_ref <= 14'h083b; // 'd2107
      10'd19   : out_data_ref <= 14'h07fc; // 'd2044
      10'd20   : out_data_ref <= 14'h0480; // 'd1152
      10'd21   : out_data_ref <= 14'h0065; // 'd101
      10'd22   : out_data_ref <= 14'h0d6f; // 'd3439
      10'd23   : out_data_ref <= 14'h0700; // 'd1792
      10'd24   : out_data_ref <= 14'h0f21; // 'd3873
      10'd25   : out_data_ref <= 14'h0d2c; // 'd3372
      10'd26   : out_data_ref <= 14'h00f6; // 'd246
      10'd27   : out_data_ref <= 14'h0363; // 'd867
      10'd28   : out_data_ref <= 14'h005b; // 'd91
      10'd29   : out_data_ref <= 14'h02fb; // 'd763
      10'd30   : out_data_ref <= 14'h0cee; // 'd3310
      10'd31   : out_data_ref <= 14'h10ea; // 'd4330
      10'd32   : out_data_ref <= 14'h07ac; // 'd1964
      10'd33   : out_data_ref <= 14'h043b; // 'd1083
      10'd34   : out_data_ref <= 14'h0993; // 'd2451
      10'd35   : out_data_ref <= 14'h0751; // 'd1873
      10'd36   : out_data_ref <= 14'h004c; // 'd76
      10'd37   : out_data_ref <= 14'h0097; // 'd151
      10'd38   : out_data_ref <= 14'h0225; // 'd549
      10'd39   : out_data_ref <= 14'h0686; // 'd1670
      10'd40   : out_data_ref <= 14'h0ee9; // 'd3817
      10'd41   : out_data_ref <= 14'h0582; // 'd1410
      10'd42   : out_data_ref <= 14'h0005; // 'd5
      10'd43   : out_data_ref <= 14'h052e; // 'd1326
      10'd44   : out_data_ref <= 14'h0adf; // 'd2783
      10'd45   : out_data_ref <= 14'h109e; // 'd4254
      10'd46   : out_data_ref <= 14'h0cd9; // 'd3289
      10'd47   : out_data_ref <= 14'h11b8; // 'd4536
      10'd48   : out_data_ref <= 14'h0fc0; // 'd4032
      10'd49   : out_data_ref <= 14'h0abe; // 'd2750
      10'd50   : out_data_ref <= 14'h0bf0; // 'd3056
      10'd51   : out_data_ref <= 14'h0500; // 'd1280
      10'd52   : out_data_ref <= 14'h07cc; // 'd1996
      10'd53   : out_data_ref <= 14'h0d0b; // 'd3339
      10'd54   : out_data_ref <= 14'h024b; // 'd587
      10'd55   : out_data_ref <= 14'h06ce; // 'd1742
      10'd56   : out_data_ref <= 14'h0255; // 'd597
      10'd57   : out_data_ref <= 14'h0d08; // 'd3336
      10'd58   : out_data_ref <= 14'h099e; // 'd2462
      10'd59   : out_data_ref <= 14'h0ce3; // 'd3299
      10'd60   : out_data_ref <= 14'h05bd; // 'd1469
      10'd61   : out_data_ref <= 14'h0b48; // 'd2888
      10'd62   : out_data_ref <= 14'h0fbb; // 'd4027
      10'd63   : out_data_ref <= 14'h0895; // 'd2197
      10'd64   : out_data_ref <= 14'h09ae; // 'd2478
      10'd65   : out_data_ref <= 14'h07ec; // 'd2028
      10'd66   : out_data_ref <= 14'h090e; // 'd2318
      10'd67   : out_data_ref <= 14'h00eb; // 'd235
      10'd68   : out_data_ref <= 14'h086e; // 'd2158
      10'd69   : out_data_ref <= 14'h097c; // 'd2428
      10'd70   : out_data_ref <= 14'h063f; // 'd1599
      10'd71   : out_data_ref <= 14'h0593; // 'd1427
      10'd72   : out_data_ref <= 14'h026f; // 'd623
      10'd73   : out_data_ref <= 14'h02de; // 'd734
      10'd74   : out_data_ref <= 14'h112a; // 'd4394
      10'd75   : out_data_ref <= 14'h103e; // 'd4158
      10'd76   : out_data_ref <= 14'h0097; // 'd151
      10'd77   : out_data_ref <= 14'h04c1; // 'd1217
      10'd78   : out_data_ref <= 14'h03d4; // 'd980
      10'd79   : out_data_ref <= 14'h0e5c; // 'd3676
      10'd80   : out_data_ref <= 14'h0532; // 'd1330
      10'd81   : out_data_ref <= 14'h0469; // 'd1129
      10'd82   : out_data_ref <= 14'h0b5c; // 'd2908
      10'd83   : out_data_ref <= 14'h00ff; // 'd255
      10'd84   : out_data_ref <= 14'h1153; // 'd4435
      10'd85   : out_data_ref <= 14'h0f1b; // 'd3867
      10'd86   : out_data_ref <= 14'h0500; // 'd1280
      10'd87   : out_data_ref <= 14'h0b1b; // 'd2843
      10'd88   : out_data_ref <= 14'h049e; // 'd1182
      10'd89   : out_data_ref <= 14'h06c7; // 'd1735
      10'd90   : out_data_ref <= 14'h0603; // 'd1539
      10'd91   : out_data_ref <= 14'h1148; // 'd4424
      10'd92   : out_data_ref <= 14'h102e; // 'd4142
      10'd93   : out_data_ref <= 14'h0ed1; // 'd3793
      10'd94   : out_data_ref <= 14'h085e; // 'd2142
      10'd95   : out_data_ref <= 14'h084c; // 'd2124
      10'd96   : out_data_ref <= 14'h052f; // 'd1327
      10'd97   : out_data_ref <= 14'h0f7b; // 'd3963
      10'd98   : out_data_ref <= 14'h0f20; // 'd3872
      10'd99   : out_data_ref <= 14'h06ad; // 'd1709
      10'd100  : out_data_ref <= 14'h0a2a; // 'd2602
      10'd101  : out_data_ref <= 14'h0482; // 'd1154
      10'd102  : out_data_ref <= 14'h057d; // 'd1405
      10'd103  : out_data_ref <= 14'h04de; // 'd1246
      10'd104  : out_data_ref <= 14'h06ef; // 'd1775
      10'd105  : out_data_ref <= 14'h0abc; // 'd2748
      10'd106  : out_data_ref <= 14'h08fe; // 'd2302
      10'd107  : out_data_ref <= 14'h0674; // 'd1652
      10'd108  : out_data_ref <= 14'h0e8b; // 'd3723
      10'd109  : out_data_ref <= 14'h0e26; // 'd3622
      10'd110  : out_data_ref <= 14'h02f7; // 'd759
      10'd111  : out_data_ref <= 14'h1152; // 'd4434
      10'd112  : out_data_ref <= 14'h017a; // 'd378
      10'd113  : out_data_ref <= 14'h0406; // 'd1030
      10'd114  : out_data_ref <= 14'h0cc1; // 'd3265
      10'd115  : out_data_ref <= 14'h0220; // 'd544
      10'd116  : out_data_ref <= 14'h067e; // 'd1662
      10'd117  : out_data_ref <= 14'h0917; // 'd2327
      10'd118  : out_data_ref <= 14'h11c0; // 'd4544
      10'd119  : out_data_ref <= 14'h0d8f; // 'd3471
      10'd120  : out_data_ref <= 14'h112b; // 'd4395
      10'd121  : out_data_ref <= 14'h0c67; // 'd3175
      10'd122  : out_data_ref <= 14'h06ce; // 'd1742
      10'd123  : out_data_ref <= 14'h0016; // 'd22
      10'd124  : out_data_ref <= 14'h00ad; // 'd173
      10'd125  : out_data_ref <= 14'h0d19; // 'd3353
      10'd126  : out_data_ref <= 14'h01d6; // 'd470
      10'd127  : out_data_ref <= 14'h0b49; // 'd2889
      10'd128  : out_data_ref <= 14'h1158; // 'd4440
      10'd129  : out_data_ref <= 14'h0e95; // 'd3733
      10'd130  : out_data_ref <= 14'h0abd; // 'd2749
      10'd131  : out_data_ref <= 14'h11c5; // 'd4549
      10'd132  : out_data_ref <= 14'h0e3d; // 'd3645
      10'd133  : out_data_ref <= 14'h0dcc; // 'd3532
      10'd134  : out_data_ref <= 14'h0e30; // 'd3632
      10'd135  : out_data_ref <= 14'h0f93; // 'd3987
      10'd136  : out_data_ref <= 14'h10fa; // 'd4346
      10'd137  : out_data_ref <= 14'h0f29; // 'd3881
      10'd138  : out_data_ref <= 14'h0627; // 'd1575
      10'd139  : out_data_ref <= 14'h1168; // 'd4456
      10'd140  : out_data_ref <= 14'h0b70; // 'd2928
      10'd141  : out_data_ref <= 14'h0d5b; // 'd3419
      10'd142  : out_data_ref <= 14'h0d7c; // 'd3452
      10'd143  : out_data_ref <= 14'h0370; // 'd880
      10'd144  : out_data_ref <= 14'h04c1; // 'd1217
      10'd145  : out_data_ref <= 14'h02e1; // 'd737
      10'd146  : out_data_ref <= 14'h0cbf; // 'd3263
      10'd147  : out_data_ref <= 14'h0bf0; // 'd3056
      10'd148  : out_data_ref <= 14'h0901; // 'd2305
      10'd149  : out_data_ref <= 14'h0a8c; // 'd2700
      10'd150  : out_data_ref <= 14'h052c; // 'd1324
      10'd151  : out_data_ref <= 14'h06aa; // 'd1706
      10'd152  : out_data_ref <= 14'h0e51; // 'd3665
      10'd153  : out_data_ref <= 14'h1201; // 'd4609
      10'd154  : out_data_ref <= 14'h0b40; // 'd2880
      10'd155  : out_data_ref <= 14'h0f5a; // 'd3930
      10'd156  : out_data_ref <= 14'h0161; // 'd353
      10'd157  : out_data_ref <= 14'h0aa3; // 'd2723
      10'd158  : out_data_ref <= 14'h0851; // 'd2129
      10'd159  : out_data_ref <= 14'h065e; // 'd1630
      10'd160  : out_data_ref <= 14'h0f0c; // 'd3852
      10'd161  : out_data_ref <= 14'h0d4a; // 'd3402
      10'd162  : out_data_ref <= 14'h0ed4; // 'd3796
      10'd163  : out_data_ref <= 14'h1115; // 'd4373
      10'd164  : out_data_ref <= 14'h027a; // 'd634
      10'd165  : out_data_ref <= 14'h105b; // 'd4187
      10'd166  : out_data_ref <= 14'h0032; // 'd50
      10'd167  : out_data_ref <= 14'h0f69; // 'd3945
      10'd168  : out_data_ref <= 14'h0a66; // 'd2662
      10'd169  : out_data_ref <= 14'h0804; // 'd2052
      10'd170  : out_data_ref <= 14'h08f4; // 'd2292
      10'd171  : out_data_ref <= 14'h10c3; // 'd4291
      10'd172  : out_data_ref <= 14'h0001; // 'd1
      10'd173  : out_data_ref <= 14'h0eba; // 'd3770
      10'd174  : out_data_ref <= 14'h07d9; // 'd2009
      10'd175  : out_data_ref <= 14'h0050; // 'd80
      10'd176  : out_data_ref <= 14'h106e; // 'd4206
      10'd177  : out_data_ref <= 14'h0fca; // 'd4042
      10'd178  : out_data_ref <= 14'h00b5; // 'd181
      10'd179  : out_data_ref <= 14'h04c3; // 'd1219
      10'd180  : out_data_ref <= 14'h1137; // 'd4407
      10'd181  : out_data_ref <= 14'h104c; // 'd4172
      10'd182  : out_data_ref <= 14'h0a37; // 'd2615
      10'd183  : out_data_ref <= 14'h0c4b; // 'd3147
      10'd184  : out_data_ref <= 14'h02d6; // 'd726
      10'd185  : out_data_ref <= 14'h0414; // 'd1044
      10'd186  : out_data_ref <= 14'h0cd6; // 'd3286
      10'd187  : out_data_ref <= 14'h0118; // 'd280
      10'd188  : out_data_ref <= 14'h04b5; // 'd1205
      10'd189  : out_data_ref <= 14'h11e6; // 'd4582
      10'd190  : out_data_ref <= 14'h0227; // 'd551
      10'd191  : out_data_ref <= 14'h0d83; // 'd3459
      10'd192  : out_data_ref <= 14'h0524; // 'd1316
      10'd193  : out_data_ref <= 14'h10ba; // 'd4282
      10'd194  : out_data_ref <= 14'h023f; // 'd575
      10'd195  : out_data_ref <= 14'h10c0; // 'd4288
      10'd196  : out_data_ref <= 14'h0a09; // 'd2569
      10'd197  : out_data_ref <= 14'h016c; // 'd364
      10'd198  : out_data_ref <= 14'h011e; // 'd286
      10'd199  : out_data_ref <= 14'h0ca8; // 'd3240
      10'd200  : out_data_ref <= 14'h0c48; // 'd3144
      10'd201  : out_data_ref <= 14'h018a; // 'd394
      10'd202  : out_data_ref <= 14'h017e; // 'd382
      10'd203  : out_data_ref <= 14'h07b7; // 'd1975
      10'd204  : out_data_ref <= 14'h0f5c; // 'd3932
      10'd205  : out_data_ref <= 14'h0b12; // 'd2834
      10'd206  : out_data_ref <= 14'h0e53; // 'd3667
      10'd207  : out_data_ref <= 14'h109a; // 'd4250
      10'd208  : out_data_ref <= 14'h04f4; // 'd1268
      10'd209  : out_data_ref <= 14'h0477; // 'd1143
      10'd210  : out_data_ref <= 14'h09cd; // 'd2509
      10'd211  : out_data_ref <= 14'h09ec; // 'd2540
      10'd212  : out_data_ref <= 14'h01fb; // 'd507
      10'd213  : out_data_ref <= 14'h0c07; // 'd3079
      10'd214  : out_data_ref <= 14'h0faa; // 'd4010
      10'd215  : out_data_ref <= 14'h09de; // 'd2526
      10'd216  : out_data_ref <= 14'h0932; // 'd2354
      10'd217  : out_data_ref <= 14'h0690; // 'd1680
      10'd218  : out_data_ref <= 14'h04a8; // 'd1192
      10'd219  : out_data_ref <= 14'h0b0a; // 'd2826
      10'd220  : out_data_ref <= 14'h0b4d; // 'd2893
      10'd221  : out_data_ref <= 14'h00b5; // 'd181
      10'd222  : out_data_ref <= 14'h033a; // 'd826
      10'd223  : out_data_ref <= 14'h07f0; // 'd2032
      10'd224  : out_data_ref <= 14'h0171; // 'd369
      10'd225  : out_data_ref <= 14'h0208; // 'd520
      10'd226  : out_data_ref <= 14'h0ee2; // 'd3810
      10'd227  : out_data_ref <= 14'h0687; // 'd1671
      10'd228  : out_data_ref <= 14'h06ae; // 'd1710
      10'd229  : out_data_ref <= 14'h0652; // 'd1618
      10'd230  : out_data_ref <= 14'h093a; // 'd2362
      10'd231  : out_data_ref <= 14'h0fc3; // 'd4035
      10'd232  : out_data_ref <= 14'h0a7e; // 'd2686
      10'd233  : out_data_ref <= 14'h0df3; // 'd3571
      10'd234  : out_data_ref <= 14'h06f8; // 'd1784
      10'd235  : out_data_ref <= 14'h00da; // 'd218
      10'd236  : out_data_ref <= 14'h0803; // 'd2051
      10'd237  : out_data_ref <= 14'h0e49; // 'd3657
      10'd238  : out_data_ref <= 14'h0a3b; // 'd2619
      10'd239  : out_data_ref <= 14'h0d70; // 'd3440
      10'd240  : out_data_ref <= 14'h0d87; // 'd3463
      10'd241  : out_data_ref <= 14'h064d; // 'd1613
      10'd242  : out_data_ref <= 14'h020f; // 'd527
      10'd243  : out_data_ref <= 14'h0fc3; // 'd4035
      10'd244  : out_data_ref <= 14'h0534; // 'd1332
      10'd245  : out_data_ref <= 14'h11ef; // 'd4591
      10'd246  : out_data_ref <= 14'h114f; // 'd4431
      10'd247  : out_data_ref <= 14'h0b7a; // 'd2938
      10'd248  : out_data_ref <= 14'h0204; // 'd516
      10'd249  : out_data_ref <= 14'h0b8d; // 'd2957
      10'd250  : out_data_ref <= 14'h0bba; // 'd3002
      10'd251  : out_data_ref <= 14'h0dd4; // 'd3540
      10'd252  : out_data_ref <= 14'h0d7a; // 'd3450
      10'd253  : out_data_ref <= 14'h0006; // 'd6
      10'd254  : out_data_ref <= 14'h052c; // 'd1324
      10'd255  : out_data_ref <= 14'h0e79; // 'd3705
      10'd256  : out_data_ref <= 14'h03e4; // 'd996
      10'd257  : out_data_ref <= 14'h055d; // 'd1373
      10'd258  : out_data_ref <= 14'h0125; // 'd293
      10'd259  : out_data_ref <= 14'h066b; // 'd1643
      10'd260  : out_data_ref <= 14'h0d79; // 'd3449
      10'd261  : out_data_ref <= 14'h04f9; // 'd1273
      10'd262  : out_data_ref <= 14'h066f; // 'd1647
      10'd263  : out_data_ref <= 14'h038a; // 'd906
      10'd264  : out_data_ref <= 14'h0a12; // 'd2578
      10'd265  : out_data_ref <= 14'h08f8; // 'd2296
      10'd266  : out_data_ref <= 14'h043d; // 'd1085
      10'd267  : out_data_ref <= 14'h0dc2; // 'd3522
      10'd268  : out_data_ref <= 14'h0089; // 'd137
      10'd269  : out_data_ref <= 14'h031a; // 'd794
      10'd270  : out_data_ref <= 14'h078e; // 'd1934
      10'd271  : out_data_ref <= 14'h0886; // 'd2182
      10'd272  : out_data_ref <= 14'h1016; // 'd4118
      10'd273  : out_data_ref <= 14'h016e; // 'd366
      10'd274  : out_data_ref <= 14'h0031; // 'd49
      10'd275  : out_data_ref <= 14'h0725; // 'd1829
      10'd276  : out_data_ref <= 14'h0a01; // 'd2561
      10'd277  : out_data_ref <= 14'h03f7; // 'd1015
      10'd278  : out_data_ref <= 14'h01c2; // 'd450
      10'd279  : out_data_ref <= 14'h06c0; // 'd1728
      10'd280  : out_data_ref <= 14'h0bc7; // 'd3015
      10'd281  : out_data_ref <= 14'h0c96; // 'd3222
      10'd282  : out_data_ref <= 14'h0cce; // 'd3278
      10'd283  : out_data_ref <= 14'h10ad; // 'd4269
      10'd284  : out_data_ref <= 14'h085e; // 'd2142
      10'd285  : out_data_ref <= 14'h0ff9; // 'd4089
      10'd286  : out_data_ref <= 14'h0968; // 'd2408
      10'd287  : out_data_ref <= 14'h0797; // 'd1943
      10'd288  : out_data_ref <= 14'h11c8; // 'd4552
      10'd289  : out_data_ref <= 14'h0a69; // 'd2665
      10'd290  : out_data_ref <= 14'h01de; // 'd478
      10'd291  : out_data_ref <= 14'h0e63; // 'd3683
      10'd292  : out_data_ref <= 14'h04c8; // 'd1224
      10'd293  : out_data_ref <= 14'h0a3c; // 'd2620
      10'd294  : out_data_ref <= 14'h0d1a; // 'd3354
      10'd295  : out_data_ref <= 14'h0f1c; // 'd3868
      10'd296  : out_data_ref <= 14'h0edd; // 'd3805
      10'd297  : out_data_ref <= 14'h03dc; // 'd988
      10'd298  : out_data_ref <= 14'h0550; // 'd1360
      10'd299  : out_data_ref <= 14'h0e91; // 'd3729
      10'd300  : out_data_ref <= 14'h0d64; // 'd3428
      10'd301  : out_data_ref <= 14'h1133; // 'd4403
      10'd302  : out_data_ref <= 14'h00c8; // 'd200
      10'd303  : out_data_ref <= 14'h09df; // 'd2527
      10'd304  : out_data_ref <= 14'h04fb; // 'd1275
      10'd305  : out_data_ref <= 14'h1183; // 'd4483
      10'd306  : out_data_ref <= 14'h06b2; // 'd1714
      10'd307  : out_data_ref <= 14'h05c6; // 'd1478
      10'd308  : out_data_ref <= 14'h0150; // 'd336
      10'd309  : out_data_ref <= 14'h0bf1; // 'd3057
      10'd310  : out_data_ref <= 14'h03e0; // 'd992
      10'd311  : out_data_ref <= 14'h088d; // 'd2189
      10'd312  : out_data_ref <= 14'h061a; // 'd1562
      10'd313  : out_data_ref <= 14'h0a06; // 'd2566
      10'd314  : out_data_ref <= 14'h0ba1; // 'd2977
      10'd315  : out_data_ref <= 14'h0817; // 'd2071
      10'd316  : out_data_ref <= 14'h03c7; // 'd967
      10'd317  : out_data_ref <= 14'h1163; // 'd4451
      10'd318  : out_data_ref <= 14'h063a; // 'd1594
      10'd319  : out_data_ref <= 14'h0c83; // 'd3203
      10'd320  : out_data_ref <= 14'h0373; // 'd883
      10'd321  : out_data_ref <= 14'h05c5; // 'd1477
      10'd322  : out_data_ref <= 14'h009c; // 'd156
      10'd323  : out_data_ref <= 14'h119e; // 'd4510
      10'd324  : out_data_ref <= 14'h0a8c; // 'd2700
      10'd325  : out_data_ref <= 14'h0bb4; // 'd2996
      10'd326  : out_data_ref <= 14'h0c86; // 'd3206
      10'd327  : out_data_ref <= 14'h0c8b; // 'd3211
      10'd328  : out_data_ref <= 14'h0fa9; // 'd4009
      10'd329  : out_data_ref <= 14'h0a29; // 'd2601
      10'd330  : out_data_ref <= 14'h10b2; // 'd4274
      10'd331  : out_data_ref <= 14'h0f87; // 'd3975
      10'd332  : out_data_ref <= 14'h0333; // 'd819
      10'd333  : out_data_ref <= 14'h03c5; // 'd965
      10'd334  : out_data_ref <= 14'h074a; // 'd1866
      10'd335  : out_data_ref <= 14'h088d; // 'd2189
      10'd336  : out_data_ref <= 14'h0ca9; // 'd3241
      10'd337  : out_data_ref <= 14'h0bcf; // 'd3023
      10'd338  : out_data_ref <= 14'h0716; // 'd1814
      10'd339  : out_data_ref <= 14'h0a55; // 'd2645
      10'd340  : out_data_ref <= 14'h0933; // 'd2355
      10'd341  : out_data_ref <= 14'h0853; // 'd2131
      10'd342  : out_data_ref <= 14'h10c3; // 'd4291
      10'd343  : out_data_ref <= 14'h0d69; // 'd3433
      10'd344  : out_data_ref <= 14'h0ed7; // 'd3799
      10'd345  : out_data_ref <= 14'h0049; // 'd73
      10'd346  : out_data_ref <= 14'h0c90; // 'd3216
      10'd347  : out_data_ref <= 14'h109f; // 'd4255
      10'd348  : out_data_ref <= 14'h0ef7; // 'd3831
      10'd349  : out_data_ref <= 14'h03ce; // 'd974
      10'd350  : out_data_ref <= 14'h0c23; // 'd3107
      10'd351  : out_data_ref <= 14'h11f9; // 'd4601
      10'd352  : out_data_ref <= 14'h0798; // 'd1944
      10'd353  : out_data_ref <= 14'h0d6c; // 'd3436
      10'd354  : out_data_ref <= 14'h0efe; // 'd3838
      10'd355  : out_data_ref <= 14'h097c; // 'd2428
      10'd356  : out_data_ref <= 14'h0a33; // 'd2611
      10'd357  : out_data_ref <= 14'h00f5; // 'd245
      10'd358  : out_data_ref <= 14'h0f3d; // 'd3901
      10'd359  : out_data_ref <= 14'h0ee8; // 'd3816
      10'd360  : out_data_ref <= 14'h06fd; // 'd1789
      10'd361  : out_data_ref <= 14'h0b80; // 'd2944
      10'd362  : out_data_ref <= 14'h02a8; // 'd680
      10'd363  : out_data_ref <= 14'h1148; // 'd4424
      10'd364  : out_data_ref <= 14'h01c6; // 'd454
      10'd365  : out_data_ref <= 14'h0523; // 'd1315
      10'd366  : out_data_ref <= 14'h098a; // 'd2442
      10'd367  : out_data_ref <= 14'h0730; // 'd1840
      10'd368  : out_data_ref <= 14'h1102; // 'd4354
      10'd369  : out_data_ref <= 14'h0c19; // 'd3097
      10'd370  : out_data_ref <= 14'h008e; // 'd142
      10'd371  : out_data_ref <= 14'h05cf; // 'd1487
      10'd372  : out_data_ref <= 14'h0035; // 'd53
      10'd373  : out_data_ref <= 14'h0239; // 'd569
      10'd374  : out_data_ref <= 14'h07b8; // 'd1976
      10'd375  : out_data_ref <= 14'h098b; // 'd2443
      10'd376  : out_data_ref <= 14'h0d30; // 'd3376
      10'd377  : out_data_ref <= 14'h034a; // 'd842
      10'd378  : out_data_ref <= 14'h06c8; // 'd1736
      10'd379  : out_data_ref <= 14'h0f34; // 'd3892
      10'd380  : out_data_ref <= 14'h0e4a; // 'd3658
      10'd381  : out_data_ref <= 14'h073f; // 'd1855
      10'd382  : out_data_ref <= 14'h0153; // 'd339
      10'd383  : out_data_ref <= 14'h11bc; // 'd4540
      10'd384  : out_data_ref <= 14'h1178; // 'd4472
      10'd385  : out_data_ref <= 14'h10be; // 'd4286
      10'd386  : out_data_ref <= 14'h09c3; // 'd2499
      10'd387  : out_data_ref <= 14'h0654; // 'd1620
      10'd388  : out_data_ref <= 14'h0b33; // 'd2867
      10'd389  : out_data_ref <= 14'h0173; // 'd371
      10'd390  : out_data_ref <= 14'h059f; // 'd1439
      10'd391  : out_data_ref <= 14'h05ef; // 'd1519
      10'd392  : out_data_ref <= 14'h02fe; // 'd766
      10'd393  : out_data_ref <= 14'h0668; // 'd1640
      10'd394  : out_data_ref <= 14'h0368; // 'd872
      10'd395  : out_data_ref <= 14'h115c; // 'd4444
      10'd396  : out_data_ref <= 14'h0a31; // 'd2609
      10'd397  : out_data_ref <= 14'h003b; // 'd59
      10'd398  : out_data_ref <= 14'h0a0a; // 'd2570
      10'd399  : out_data_ref <= 14'h098e; // 'd2446
      10'd400  : out_data_ref <= 14'h08f4; // 'd2292
      10'd401  : out_data_ref <= 14'h0b16; // 'd2838
      10'd402  : out_data_ref <= 14'h0541; // 'd1345
      10'd403  : out_data_ref <= 14'h0fc6; // 'd4038
      10'd404  : out_data_ref <= 14'h03ad; // 'd941
      10'd405  : out_data_ref <= 14'h0641; // 'd1601
      10'd406  : out_data_ref <= 14'h0d52; // 'd3410
      10'd407  : out_data_ref <= 14'h021a; // 'd538
      10'd408  : out_data_ref <= 14'h0716; // 'd1814
      10'd409  : out_data_ref <= 14'h0e9b; // 'd3739
      10'd410  : out_data_ref <= 14'h0618; // 'd1560
      10'd411  : out_data_ref <= 14'h0f8d; // 'd3981
      10'd412  : out_data_ref <= 14'h0102; // 'd258
      10'd413  : out_data_ref <= 14'h0bda; // 'd3034
      10'd414  : out_data_ref <= 14'h0573; // 'd1395
      10'd415  : out_data_ref <= 14'h04ad; // 'd1197
      10'd416  : out_data_ref <= 14'h0c56; // 'd3158
      10'd417  : out_data_ref <= 14'h097c; // 'd2428
      10'd418  : out_data_ref <= 14'h08b4; // 'd2228
      10'd419  : out_data_ref <= 14'h0932; // 'd2354
      10'd420  : out_data_ref <= 14'h1048; // 'd4168
      10'd421  : out_data_ref <= 14'h0b0a; // 'd2826
      10'd422  : out_data_ref <= 14'h0064; // 'd100
      10'd423  : out_data_ref <= 14'h0805; // 'd2053
      10'd424  : out_data_ref <= 14'h0e14; // 'd3604
      10'd425  : out_data_ref <= 14'h046e; // 'd1134
      10'd426  : out_data_ref <= 14'h0adb; // 'd2779
      10'd427  : out_data_ref <= 14'h019c; // 'd412
      10'd428  : out_data_ref <= 14'h0d1d; // 'd3357
      10'd429  : out_data_ref <= 14'h0dcf; // 'd3535
      10'd430  : out_data_ref <= 14'h1090; // 'd4240
      10'd431  : out_data_ref <= 14'h0f8a; // 'd3978
      10'd432  : out_data_ref <= 14'h0f09; // 'd3849
      10'd433  : out_data_ref <= 14'h04a4; // 'd1188
      10'd434  : out_data_ref <= 14'h0565; // 'd1381
      10'd435  : out_data_ref <= 14'h06a1; // 'd1697
      10'd436  : out_data_ref <= 14'h0af8; // 'd2808
      10'd437  : out_data_ref <= 14'h014f; // 'd335
      10'd438  : out_data_ref <= 14'h0ba5; // 'd2981
      10'd439  : out_data_ref <= 14'h0d6c; // 'd3436
      10'd440  : out_data_ref <= 14'h0d72; // 'd3442
      10'd441  : out_data_ref <= 14'h088c; // 'd2188
      10'd442  : out_data_ref <= 14'h0f3d; // 'd3901
      10'd443  : out_data_ref <= 14'h02f3; // 'd755
      10'd444  : out_data_ref <= 14'h0a24; // 'd2596
      10'd445  : out_data_ref <= 14'h0f51; // 'd3921
      10'd446  : out_data_ref <= 14'h0f9b; // 'd3995
      10'd447  : out_data_ref <= 14'h0415; // 'd1045
      10'd448  : out_data_ref <= 14'h0b3f; // 'd2879
      10'd449  : out_data_ref <= 14'h11a9; // 'd4521
      10'd450  : out_data_ref <= 14'h07f5; // 'd2037
      10'd451  : out_data_ref <= 14'h11c8; // 'd4552
      10'd452  : out_data_ref <= 14'h0ca8; // 'd3240
      10'd453  : out_data_ref <= 14'h0327; // 'd807
      10'd454  : out_data_ref <= 14'h1064; // 'd4196
      10'd455  : out_data_ref <= 14'h06fd; // 'd1789
      10'd456  : out_data_ref <= 14'h0dc8; // 'd3528
      10'd457  : out_data_ref <= 14'h0275; // 'd629
      10'd458  : out_data_ref <= 14'h0f53; // 'd3923
      10'd459  : out_data_ref <= 14'h07f1; // 'd2033
      10'd460  : out_data_ref <= 14'h0b4e; // 'd2894
      10'd461  : out_data_ref <= 14'h07b9; // 'd1977
      10'd462  : out_data_ref <= 14'h0156; // 'd342
      10'd463  : out_data_ref <= 14'h10d4; // 'd4308
      10'd464  : out_data_ref <= 14'h0eab; // 'd3755
      10'd465  : out_data_ref <= 14'h1081; // 'd4225
      10'd466  : out_data_ref <= 14'h0478; // 'd1144
      10'd467  : out_data_ref <= 14'h021a; // 'd538
      10'd468  : out_data_ref <= 14'h009e; // 'd158
      10'd469  : out_data_ref <= 14'h057e; // 'd1406
      10'd470  : out_data_ref <= 14'h0254; // 'd596
      10'd471  : out_data_ref <= 14'h03ea; // 'd1002
      10'd472  : out_data_ref <= 14'h0610; // 'd1552
      10'd473  : out_data_ref <= 14'h1070; // 'd4208
      10'd474  : out_data_ref <= 14'h023f; // 'd575
      10'd475  : out_data_ref <= 14'h0312; // 'd786
      10'd476  : out_data_ref <= 14'h1109; // 'd4361
      10'd477  : out_data_ref <= 14'h07e8; // 'd2024
      10'd478  : out_data_ref <= 14'h0d47; // 'd3399
      10'd479  : out_data_ref <= 14'h10ca; // 'd4298
      10'd480  : out_data_ref <= 14'h0c72; // 'd3186
      10'd481  : out_data_ref <= 14'h0eed; // 'd3821
      10'd482  : out_data_ref <= 14'h0935; // 'd2357
      10'd483  : out_data_ref <= 14'h0b9d; // 'd2973
      10'd484  : out_data_ref <= 14'h0250; // 'd592
      10'd485  : out_data_ref <= 14'h056b; // 'd1387
      10'd486  : out_data_ref <= 14'h0df7; // 'd3575
      10'd487  : out_data_ref <= 14'h0a15; // 'd2581
      10'd488  : out_data_ref <= 14'h0ada; // 'd2778
      10'd489  : out_data_ref <= 14'h0b8a; // 'd2954
      10'd490  : out_data_ref <= 14'h0b85; // 'd2949
      10'd491  : out_data_ref <= 14'h0cde; // 'd3294
      10'd492  : out_data_ref <= 14'h0efc; // 'd3836
      10'd493  : out_data_ref <= 14'h0bfa; // 'd3066
      10'd494  : out_data_ref <= 14'h0bc2; // 'd3010
      10'd495  : out_data_ref <= 14'h10bf; // 'd4287
      10'd496  : out_data_ref <= 14'h01d2; // 'd466
      10'd497  : out_data_ref <= 14'h0d0b; // 'd3339
      10'd498  : out_data_ref <= 14'h0727; // 'd1831
      10'd499  : out_data_ref <= 14'h0bf8; // 'd3064
      10'd500  : out_data_ref <= 14'h0585; // 'd1413
      10'd501  : out_data_ref <= 14'h0670; // 'd1648
      10'd502  : out_data_ref <= 14'h0c94; // 'd3220
      10'd503  : out_data_ref <= 14'h0a12; // 'd2578
      10'd504  : out_data_ref <= 14'h008f; // 'd143
      10'd505  : out_data_ref <= 14'h02d7; // 'd727
      10'd506  : out_data_ref <= 14'h0dbc; // 'd3516
      10'd507  : out_data_ref <= 14'h1038; // 'd4152
      10'd508  : out_data_ref <= 14'h00a7; // 'd167
      10'd509  : out_data_ref <= 14'h040e; // 'd1038
      10'd510  : out_data_ref <= 14'h0b7d; // 'd2941
      10'd511  : out_data_ref <= 14'h0942; // 'd2370
      10'd512  : out_data_ref <= 14'h0591; // 'd1425
      10'd513  : out_data_ref <= 14'h0a5d; // 'd2653
      10'd514  : out_data_ref <= 14'h09cd; // 'd2509
      10'd515  : out_data_ref <= 14'h0f7f; // 'd3967
      10'd516  : out_data_ref <= 14'h077a; // 'd1914
      10'd517  : out_data_ref <= 14'h0ea2; // 'd3746
      10'd518  : out_data_ref <= 14'h06f0; // 'd1776
      10'd519  : out_data_ref <= 14'h102a; // 'd4138
      10'd520  : out_data_ref <= 14'h05cb; // 'd1483
      10'd521  : out_data_ref <= 14'h0c4b; // 'd3147
      10'd522  : out_data_ref <= 14'h1191; // 'd4497
      10'd523  : out_data_ref <= 14'h0279; // 'd633
      10'd524  : out_data_ref <= 14'h0d56; // 'd3414
      10'd525  : out_data_ref <= 14'h02c1; // 'd705
      10'd526  : out_data_ref <= 14'h1057; // 'd4183
      10'd527  : out_data_ref <= 14'h0e3d; // 'd3645
      10'd528  : out_data_ref <= 14'h11b9; // 'd4537
      10'd529  : out_data_ref <= 14'h0955; // 'd2389
      10'd530  : out_data_ref <= 14'h0320; // 'd800
      10'd531  : out_data_ref <= 14'h0366; // 'd870
      10'd532  : out_data_ref <= 14'h071d; // 'd1821
      10'd533  : out_data_ref <= 14'h04a9; // 'd1193
      10'd534  : out_data_ref <= 14'h105c; // 'd4188
      10'd535  : out_data_ref <= 14'h0f25; // 'd3877
      10'd536  : out_data_ref <= 14'h0693; // 'd1683
      10'd537  : out_data_ref <= 14'h0e0d; // 'd3597
      10'd538  : out_data_ref <= 14'h0f41; // 'd3905
      10'd539  : out_data_ref <= 14'h11a6; // 'd4518
      10'd540  : out_data_ref <= 14'h09d6; // 'd2518
      10'd541  : out_data_ref <= 14'h06f7; // 'd1783
      10'd542  : out_data_ref <= 14'h03ed; // 'd1005
      10'd543  : out_data_ref <= 14'h10a4; // 'd4260
      10'd544  : out_data_ref <= 14'h1038; // 'd4152
      10'd545  : out_data_ref <= 14'h1004; // 'd4100
      10'd546  : out_data_ref <= 14'h07c4; // 'd1988
      10'd547  : out_data_ref <= 14'h0c74; // 'd3188
      10'd548  : out_data_ref <= 14'h0be7; // 'd3047
      10'd549  : out_data_ref <= 14'h114f; // 'd4431
      10'd550  : out_data_ref <= 14'h0aa8; // 'd2728
      10'd551  : out_data_ref <= 14'h0414; // 'd1044
      10'd552  : out_data_ref <= 14'h05fc; // 'd1532
      10'd553  : out_data_ref <= 14'h03b6; // 'd950
      10'd554  : out_data_ref <= 14'h084c; // 'd2124
      10'd555  : out_data_ref <= 14'h02f1; // 'd753
      10'd556  : out_data_ref <= 14'h0993; // 'd2451
      10'd557  : out_data_ref <= 14'h0d2b; // 'd3371
      10'd558  : out_data_ref <= 14'h0aa2; // 'd2722
      10'd559  : out_data_ref <= 14'h09e7; // 'd2535
      10'd560  : out_data_ref <= 14'h04de; // 'd1246
      10'd561  : out_data_ref <= 14'h03c6; // 'd966
      10'd562  : out_data_ref <= 14'h1071; // 'd4209
      10'd563  : out_data_ref <= 14'h0680; // 'd1664
      10'd564  : out_data_ref <= 14'h015c; // 'd348
      10'd565  : out_data_ref <= 14'h083b; // 'd2107
      10'd566  : out_data_ref <= 14'h07fd; // 'd2045
      10'd567  : out_data_ref <= 14'h070e; // 'd1806
      10'd568  : out_data_ref <= 14'h0be4; // 'd3044
      10'd569  : out_data_ref <= 14'h0c14; // 'd3092
      10'd570  : out_data_ref <= 14'h0ba8; // 'd2984
      10'd571  : out_data_ref <= 14'h0818; // 'd2072
      10'd572  : out_data_ref <= 14'h010c; // 'd268
      10'd573  : out_data_ref <= 14'h0ffb; // 'd4091
      10'd574  : out_data_ref <= 14'h0e7c; // 'd3708
      10'd575  : out_data_ref <= 14'h0e10; // 'd3600
      10'd576  : out_data_ref <= 14'h0add; // 'd2781
      10'd577  : out_data_ref <= 14'h116a; // 'd4458
      10'd578  : out_data_ref <= 14'h0125; // 'd293
      10'd579  : out_data_ref <= 14'h069d; // 'd1693
      10'd580  : out_data_ref <= 14'h07d4; // 'd2004
      10'd581  : out_data_ref <= 14'h0777; // 'd1911
      10'd582  : out_data_ref <= 14'h0b0b; // 'd2827
      10'd583  : out_data_ref <= 14'h0f65; // 'd3941
      10'd584  : out_data_ref <= 14'h04b1; // 'd1201
      10'd585  : out_data_ref <= 14'h0a03; // 'd2563
      10'd586  : out_data_ref <= 14'h099a; // 'd2458
      10'd587  : out_data_ref <= 14'h10a2; // 'd4258
      10'd588  : out_data_ref <= 14'h0707; // 'd1799
      10'd589  : out_data_ref <= 14'h0080; // 'd128
      10'd590  : out_data_ref <= 14'h071c; // 'd1820
      10'd591  : out_data_ref <= 14'h0c04; // 'd3076
      10'd592  : out_data_ref <= 14'h1115; // 'd4373
      10'd593  : out_data_ref <= 14'h02fb; // 'd763
      10'd594  : out_data_ref <= 14'h0d69; // 'd3433
      10'd595  : out_data_ref <= 14'h09b3; // 'd2483
      10'd596  : out_data_ref <= 14'h08e8; // 'd2280
      10'd597  : out_data_ref <= 14'h09d2; // 'd2514
      10'd598  : out_data_ref <= 14'h10bc; // 'd4284
      10'd599  : out_data_ref <= 14'h0763; // 'd1891
      10'd600  : out_data_ref <= 14'h063f; // 'd1599
      10'd601  : out_data_ref <= 14'h0be7; // 'd3047
      10'd602  : out_data_ref <= 14'h0dc2; // 'd3522
      10'd603  : out_data_ref <= 14'h0ef5; // 'd3829
      10'd604  : out_data_ref <= 14'h040d; // 'd1037
      10'd605  : out_data_ref <= 14'h0a0e; // 'd2574
      10'd606  : out_data_ref <= 14'h0d4e; // 'd3406
      10'd607  : out_data_ref <= 14'h05db; // 'd1499
      10'd608  : out_data_ref <= 14'h02f5; // 'd757
      10'd609  : out_data_ref <= 14'h0406; // 'd1030
      10'd610  : out_data_ref <= 14'h1189; // 'd4489
      10'd611  : out_data_ref <= 14'h0d5b; // 'd3419
      10'd612  : out_data_ref <= 14'h119b; // 'd4507
      10'd613  : out_data_ref <= 14'h0835; // 'd2101
      10'd614  : out_data_ref <= 14'h03aa; // 'd938
      10'd615  : out_data_ref <= 14'h01d5; // 'd469
      10'd616  : out_data_ref <= 14'h01b9; // 'd441
      10'd617  : out_data_ref <= 14'h1098; // 'd4248
      10'd618  : out_data_ref <= 14'h10ec; // 'd4332
      10'd619  : out_data_ref <= 14'h00a7; // 'd167
      10'd620  : out_data_ref <= 14'h04b9; // 'd1209
      10'd621  : out_data_ref <= 14'h0109; // 'd265
      10'd622  : out_data_ref <= 14'h0e67; // 'd3687
      10'd623  : out_data_ref <= 14'h04d0; // 'd1232
      10'd624  : out_data_ref <= 14'h0645; // 'd1605
      10'd625  : out_data_ref <= 14'h094e; // 'd2382
      10'd626  : out_data_ref <= 14'h03fa; // 'd1018
      10'd627  : out_data_ref <= 14'h0c6b; // 'd3179
      10'd628  : out_data_ref <= 14'h0baa; // 'd2986
      10'd629  : out_data_ref <= 14'h0335; // 'd821
      10'd630  : out_data_ref <= 14'h0038; // 'd56
      10'd631  : out_data_ref <= 14'h00b1; // 'd177
      10'd632  : out_data_ref <= 14'h0899; // 'd2201
      10'd633  : out_data_ref <= 14'h0f2e; // 'd3886
      10'd634  : out_data_ref <= 14'h0fe1; // 'd4065
      10'd635  : out_data_ref <= 14'h041f; // 'd1055
      10'd636  : out_data_ref <= 14'h1097; // 'd4247
      10'd637  : out_data_ref <= 14'h09b1; // 'd2481
      10'd638  : out_data_ref <= 14'h08a3; // 'd2211
      10'd639  : out_data_ref <= 14'h0aa6; // 'd2726
      10'd640  : out_data_ref <= 14'h0955; // 'd2389
      10'd641  : out_data_ref <= 14'h0565; // 'd1381
      10'd642  : out_data_ref <= 14'h0cdb; // 'd3291
      10'd643  : out_data_ref <= 14'h08a3; // 'd2211
      10'd644  : out_data_ref <= 14'h02b1; // 'd689
      10'd645  : out_data_ref <= 14'h047e; // 'd1150
      10'd646  : out_data_ref <= 14'h0fa2; // 'd4002
      10'd647  : out_data_ref <= 14'h0c4a; // 'd3146
      10'd648  : out_data_ref <= 14'h0ffe; // 'd4094
      10'd649  : out_data_ref <= 14'h09d9; // 'd2521
      10'd650  : out_data_ref <= 14'h0402; // 'd1026
      10'd651  : out_data_ref <= 14'h05df; // 'd1503
      10'd652  : out_data_ref <= 14'h07f1; // 'd2033
      default: out_data_ref <= 14'h0;
    endcase
  end

endmodule
