module mod6343Svec35 (
    input       [34:0] z_in,
    output      [11:0] p0,
    output reg  [12:0] p1,
    output reg  [11:0] p2,
    output reg  [12:0] p3,
    output      [11:0] n0,
    output reg  [12:0] n1
) ;

    reg         [ 8:0] n0_mL;
    reg         [ 7:0] n0_Mm;

    assign p0 = z_in[11:0];

    always @ (*) begin
        case({ z_in[31], z_in[23], z_in[21], z_in[14] })
            4'h0: p1 = 13'd0;
            4'h1: p1 = 13'd3698;
            4'h2: p1 = 13'd3962;
            4'h3: p1 = 13'd1317;
            4'h4: p1 = 13'd3162;
            4'h5: p1 = 13'd517;
            4'h6: p1 = 13'd781;
            4'h7: p1 = 13'd4479;
            4'h8: p1 = 13'd3911;
            4'h9: p1 = 13'd1266;
            4'ha: p1 = 13'd1530;
            4'hb: p1 = 13'd5228;
            4'hc: p1 = 13'd730;
            4'hd: p1 = 13'd4428;
            4'he: p1 = 13'd4692;
            4'hf: p1 = 13'd2047;
        endcase
    end

    always @ (*) begin
        case({ z_in[34], z_in[32], z_in[15] })
            3'h0: p2 = 12'd0;
            3'h1: p2 = 12'd1053;
            3'h2: p2 = 12'd1479;
            3'h3: p2 = 12'd2532;
            3'h4: p2 = 12'd427;
            3'h5: p2 = 12'd1480;
            3'h6: p2 = 12'd1906;
            3'h7: p2 = 12'd2959;
        endcase
    end

    always @ (*) begin
        case({ z_in[22], z_in[20], z_in[18], z_in[13] })
            4'h0: p3 = 13'd0;
            4'h1: p3 = 13'd1849;
            4'h2: p3 = 13'd2081;
            4'h3: p3 = 13'd3930;
            4'h4: p3 = 13'd1981;
            4'h5: p3 = 13'd3830;
            4'h6: p3 = 13'd4062;
            4'h7: p3 = 13'd5911;
            4'h8: p3 = 13'd1581;
            4'h9: p3 = 13'd3430;
            4'ha: p3 = 13'd3662;
            4'hb: p3 = 13'd5511;
            4'hc: p3 = 13'd3562;
            4'hd: p3 = 13'd5411;
            4'he: p3 = 13'd5643;
            4'hf: p3 = 13'd1149;
        endcase
    end

    always @ (*) begin
        //case({ z_in[30], z_in[29], z_in[28], z_in[27], z_in[26], z_in[25], z_in[24] })
        //    7'h00: n0 = 12'h000;
        //    7'h01: n0 = 12'h003;
        //    7'h02: n0 = 12'h006;
        //    7'h03: n0 = 12'h009;
        //    7'h04: n0 = 12'h00c;
        //    7'h05: n0 = 12'h00f;
        //    7'h06: n0 = 12'h012;
        //    7'h07: n0 = 12'h015;
        //    7'h08: n0 = 12'h018;
        //    7'h09: n0 = 12'h01b;
        //    7'h0a: n0 = 12'h01e;
        //    7'h0b: n0 = 12'h021;
        //    7'h0c: n0 = 12'h024;
        //    7'h0d: n0 = 12'h027;
        //    7'h0e: n0 = 12'h02a;
        //    7'h0f: n0 = 12'h02d;
        //    7'h10: n0 = 12'h030;
        //    7'h11: n0 = 12'h033;
        //    7'h12: n0 = 12'h036;
        //    7'h13: n0 = 12'h039;
        //    7'h14: n0 = 12'h03c;
        //    7'h15: n0 = 12'h03f;
        //    7'h16: n0 = 12'h042;
        //    7'h17: n0 = 12'h045;
        //    7'h18: n0 = 12'h048;
        //    7'h19: n0 = 12'h04b;
        //    7'h1a: n0 = 12'h04e;
        //    7'h1b: n0 = 12'h051;
        //    7'h1c: n0 = 12'h054;
        //    7'h1d: n0 = 12'h057;
        //    7'h1e: n0 = 12'h05a;
        //    7'h1f: n0 = 12'h05d;
        //    7'h20: n0 = 12'h060;
        //    7'h21: n0 = 12'h063;
        //    7'h22: n0 = 12'h066;
        //    7'h23: n0 = 12'h069;
        //    7'h24: n0 = 12'h06c;
        //    7'h25: n0 = 12'h06f;
        //    7'h26: n0 = 12'h072;
        //    7'h27: n0 = 12'h075;
        //    7'h28: n0 = 12'h078;
        //    7'h29: n0 = 12'h07b;
        //    7'h2a: n0 = 12'h07e;
        //    7'h2b: n0 = 12'h081;
        //    7'h2c: n0 = 12'h084;
        //    7'h2d: n0 = 12'h087;
        //    7'h2e: n0 = 12'h08a;
        //    7'h2f: n0 = 12'h08d;
        //    7'h30: n0 = 12'h090;
        //    7'h31: n0 = 12'h093;
        //    7'h32: n0 = 12'h096;
        //    7'h33: n0 = 12'h099;
        //    7'h34: n0 = 12'h09c;
        //    7'h35: n0 = 12'h09f;
        //    7'h36: n0 = 12'h0a2;
        //    7'h37: n0 = 12'h0a5;
        //    7'h38: n0 = 12'h0a8;
        //    7'h39: n0 = 12'h0ab;
        //    7'h3a: n0 = 12'h0ae;
        //    7'h3b: n0 = 12'h0b1;
        //    7'h3c: n0 = 12'h0b4;
        //    7'h3d: n0 = 12'h0b7;
        //    7'h3e: n0 = 12'h0ba;
        //    7'h3f: n0 = 12'h0bd;
        //    7'h40: n0 = 12'h0c0;
        //    7'h41: n0 = 12'h0c3;
        //    7'h42: n0 = 12'h0c6;
        //    7'h43: n0 = 12'h0c9;
        //    7'h44: n0 = 12'h0cc;
        //    7'h45: n0 = 12'h0cf;
        //    7'h46: n0 = 12'h0d2;
        //    7'h47: n0 = 12'h0d5;
        //    7'h48: n0 = 12'h0d8;
        //    7'h49: n0 = 12'h0db;
        //    7'h4a: n0 = 12'h0de;
        //    7'h4b: n0 = 12'h0e1;
        //    7'h4c: n0 = 12'h0e4;
        //    7'h4d: n0 = 12'h0e7;
        //    7'h4e: n0 = 12'h0ea;
        //    7'h4f: n0 = 12'h0ed;
        //    7'h50: n0 = 12'h0f0;
        //    7'h51: n0 = 12'h0f3;
        //    7'h52: n0 = 12'h0f6;
        //    7'h53: n0 = 12'h0f9;
        //    7'h54: n0 = 12'h0fc;
        //    7'h55: n0 = 12'h0ff;
        //    7'h56: n0 = 12'h102;
        //    7'h57: n0 = 12'h105;
        //    7'h58: n0 = 12'h108;
        //    7'h59: n0 = 12'h10b;
        //    7'h5a: n0 = 12'h10e;
        //    7'h5b: n0 = 12'h111;
        //    7'h5c: n0 = 12'h114;
        //    7'h5d: n0 = 12'h117;
        //    7'h5e: n0 = 12'h11a;
        //    7'h5f: n0 = 12'h11d;
        //    7'h60: n0 = 12'h120;
        //    7'h61: n0 = 12'h123;
        //    7'h62: n0 = 12'h126;
        //    7'h63: n0 = 12'h129;
        //    7'h64: n0 = 12'h12c;
        //    7'h65: n0 = 12'h12f;
        //    7'h66: n0 = 12'h132;
        //    7'h67: n0 = 12'h135;
        //    7'h68: n0 = 12'h138;
        //    7'h69: n0 = 12'h13b;
        //    7'h6a: n0 = 12'h13e;
        //    7'h6b: n0 = 12'h141;
        //    7'h6c: n0 = 12'h144;
        //    7'h6d: n0 = 12'h147;
        //    7'h6e: n0 = 12'h14a;
        //    7'h6f: n0 = 12'h14d;
        //    7'h70: n0 = 12'h150;
        //    7'h71: n0 = 12'h153;
        //    7'h72: n0 = 12'h156;
        //    7'h73: n0 = 12'h159;
        //    7'h74: n0 = 12'h15c;
        //    7'h75: n0 = 12'h15f;
        //    7'h76: n0 = 12'h162;
        //    7'h77: n0 = 12'h165;
        //    7'h78: n0 = 12'h168;
        //    7'h79: n0 = 12'h16b;
        //    7'h7a: n0 = 12'h16e;
        //    7'h7b: n0 = 12'h171;
        //    7'h7c: n0 = 12'h174;
        //    7'h7d: n0 = 12'h177;
        //    7'h7e: n0 = 12'h17a;
        //    7'h7f: n0 = 12'h17d;
        //endcase
        n0_mL = { 1'b0, z_in[30:24], 1'b0 } + { 2'b0, z_in[30:24] };
        n0_Mm = { 1'b0, z_in[30:24] } + { 3'b0, n0_mL[8:4] };
    end
    assign n0 = { n0_Mm, n0_mL[3:0] };

    always @ (*) begin
        case({ z_in[33], z_in[19], z_in[17], z_in[16], z_in[12] })
            5'h00: n1 = 13'd0;
            5'h01: n1 = 13'd2247;
            5'h02: n1 = 13'd4237;
            5'h03: n1 = 13'd141;
            5'h04: n1 = 13'd2131;
            5'h05: n1 = 13'd4378;
            5'h06: n1 = 13'd25;
            5'h07: n1 = 13'd2272;
            5'h08: n1 = 13'd2181;
            5'h09: n1 = 13'd4428;
            5'h0a: n1 = 13'd75;
            5'h0b: n1 = 13'd2322;
            5'h0c: n1 = 13'd4312;
            5'h0d: n1 = 13'd216;
            5'h0e: n1 = 13'd2206;
            5'h0f: n1 = 13'd4453;
            5'h10: n1 = 13'd3385;
            5'h11: n1 = 13'd5632;
            5'h12: n1 = 13'd1279;
            5'h13: n1 = 13'd3526;
            5'h14: n1 = 13'd5516;
            5'h15: n1 = 13'd1420;
            5'h16: n1 = 13'd3410;
            5'h17: n1 = 13'd5657;
            5'h18: n1 = 13'd5566;
            5'h19: n1 = 13'd1470;
            5'h1a: n1 = 13'd3460;
            5'h1b: n1 = 13'd5707;
            5'h1c: n1 = 13'd1354;
            5'h1d: n1 = 13'd3601;
            5'h1e: n1 = 13'd5591;
            5'h1f: n1 = 13'd1495;
        endcase
    end

endmodule
