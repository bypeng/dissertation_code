module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd1277;
  localparam R_DEPTH = 'd11;
  localparam B_LEN = 'd2067;
  localparam B_DEPTH = 'd12;

  input              clk;
  input      [10: 0] in_addr;
  output reg [13: 0] in_data;
  input      [11: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      11'd0    : in_data <= 14'h1c6f; // 'd7279
      11'd1    : in_data <= 14'h1205; // 'd4613
      11'd2    : in_data <= 14'h0200; // 'd512
      11'd3    : in_data <= 14'h09e9; // 'd2537
      11'd4    : in_data <= 14'h03f4; // 'd1012
      11'd5    : in_data <= 14'h13dc; // 'd5084
      11'd6    : in_data <= 14'h1195; // 'd4501
      11'd7    : in_data <= 14'h0acf; // 'd2767
      11'd8    : in_data <= 14'h14f8; // 'd5368
      11'd9    : in_data <= 14'h1b69; // 'd7017
      11'd10   : in_data <= 14'h0b96; // 'd2966
      11'd11   : in_data <= 14'h1daf; // 'd7599
      11'd12   : in_data <= 14'h0d2a; // 'd3370
      11'd13   : in_data <= 14'h122c; // 'd4652
      11'd14   : in_data <= 14'h0025; // 'd37
      11'd15   : in_data <= 14'h061b; // 'd1563
      11'd16   : in_data <= 14'h1d8b; // 'd7563
      11'd17   : in_data <= 14'h03bb; // 'd955
      11'd18   : in_data <= 14'h048f; // 'd1167
      11'd19   : in_data <= 14'h1439; // 'd5177
      11'd20   : in_data <= 14'h11c9; // 'd4553
      11'd21   : in_data <= 14'h0e54; // 'd3668
      11'd22   : in_data <= 14'h171e; // 'd5918
      11'd23   : in_data <= 14'h0529; // 'd1321
      11'd24   : in_data <= 14'h1247; // 'd4679
      11'd25   : in_data <= 14'h1ac3; // 'd6851
      11'd26   : in_data <= 14'h1284; // 'd4740
      11'd27   : in_data <= 14'h0473; // 'd1139
      11'd28   : in_data <= 14'h10bd; // 'd4285
      11'd29   : in_data <= 14'h1011; // 'd4113
      11'd30   : in_data <= 14'h0d43; // 'd3395
      11'd31   : in_data <= 14'h1c35; // 'd7221
      11'd32   : in_data <= 14'h1e48; // 'd7752
      11'd33   : in_data <= 14'h1ced; // 'd7405
      11'd34   : in_data <= 14'h02a1; // 'd673
      11'd35   : in_data <= 14'h025f; // 'd607
      11'd36   : in_data <= 14'h172d; // 'd5933
      11'd37   : in_data <= 14'h0d32; // 'd3378
      11'd38   : in_data <= 14'h054a; // 'd1354
      11'd39   : in_data <= 14'h00bb; // 'd187
      11'd40   : in_data <= 14'h0b21; // 'd2849
      11'd41   : in_data <= 14'h1349; // 'd4937
      11'd42   : in_data <= 14'h1423; // 'd5155
      11'd43   : in_data <= 14'h1401; // 'd5121
      11'd44   : in_data <= 14'h1204; // 'd4612
      11'd45   : in_data <= 14'h0333; // 'd819
      11'd46   : in_data <= 14'h1bbd; // 'd7101
      11'd47   : in_data <= 14'h0b97; // 'd2967
      11'd48   : in_data <= 14'h0f1f; // 'd3871
      11'd49   : in_data <= 14'h09f9; // 'd2553
      11'd50   : in_data <= 14'h06d2; // 'd1746
      11'd51   : in_data <= 14'h0545; // 'd1349
      11'd52   : in_data <= 14'h1b56; // 'd6998
      11'd53   : in_data <= 14'h146b; // 'd5227
      11'd54   : in_data <= 14'h00fe; // 'd254
      11'd55   : in_data <= 14'h0fed; // 'd4077
      11'd56   : in_data <= 14'h015f; // 'd351
      11'd57   : in_data <= 14'h0ae2; // 'd2786
      11'd58   : in_data <= 14'h0605; // 'd1541
      11'd59   : in_data <= 14'h0be8; // 'd3048
      11'd60   : in_data <= 14'h1657; // 'd5719
      11'd61   : in_data <= 14'h082c; // 'd2092
      11'd62   : in_data <= 14'h03e0; // 'd992
      11'd63   : in_data <= 14'h1b0f; // 'd6927
      11'd64   : in_data <= 14'h1e65; // 'd7781
      11'd65   : in_data <= 14'h0840; // 'd2112
      11'd66   : in_data <= 14'h1ab8; // 'd6840
      11'd67   : in_data <= 14'h0dd5; // 'd3541
      11'd68   : in_data <= 14'h1805; // 'd6149
      11'd69   : in_data <= 14'h15e3; // 'd5603
      11'd70   : in_data <= 14'h0a30; // 'd2608
      11'd71   : in_data <= 14'h0ca2; // 'd3234
      11'd72   : in_data <= 14'h02be; // 'd702
      11'd73   : in_data <= 14'h10e0; // 'd4320
      11'd74   : in_data <= 14'h19a5; // 'd6565
      11'd75   : in_data <= 14'h1602; // 'd5634
      11'd76   : in_data <= 14'h1bd4; // 'd7124
      11'd77   : in_data <= 14'h054e; // 'd1358
      11'd78   : in_data <= 14'h078e; // 'd1934
      11'd79   : in_data <= 14'h19c2; // 'd6594
      11'd80   : in_data <= 14'h10d8; // 'd4312
      11'd81   : in_data <= 14'h140e; // 'd5134
      11'd82   : in_data <= 14'h0f9b; // 'd3995
      11'd83   : in_data <= 14'h1845; // 'd6213
      11'd84   : in_data <= 14'h1872; // 'd6258
      11'd85   : in_data <= 14'h12f1; // 'd4849
      11'd86   : in_data <= 14'h072b; // 'd1835
      11'd87   : in_data <= 14'h06e8; // 'd1768
      11'd88   : in_data <= 14'h0d24; // 'd3364
      11'd89   : in_data <= 14'h1dcf; // 'd7631
      11'd90   : in_data <= 14'h167d; // 'd5757
      11'd91   : in_data <= 14'h16d3; // 'd5843
      11'd92   : in_data <= 14'h0376; // 'd886
      11'd93   : in_data <= 14'h1788; // 'd6024
      11'd94   : in_data <= 14'h0f0c; // 'd3852
      11'd95   : in_data <= 14'h176d; // 'd5997
      11'd96   : in_data <= 14'h09da; // 'd2522
      11'd97   : in_data <= 14'h0033; // 'd51
      11'd98   : in_data <= 14'h0a9a; // 'd2714
      11'd99   : in_data <= 14'h13ab; // 'd5035
      11'd100  : in_data <= 14'h19ea; // 'd6634
      11'd101  : in_data <= 14'h02cf; // 'd719
      11'd102  : in_data <= 14'h1248; // 'd4680
      11'd103  : in_data <= 14'h0c98; // 'd3224
      11'd104  : in_data <= 14'h0cb8; // 'd3256
      11'd105  : in_data <= 14'h1cde; // 'd7390
      11'd106  : in_data <= 14'h0446; // 'd1094
      11'd107  : in_data <= 14'h0320; // 'd800
      11'd108  : in_data <= 14'h1e04; // 'd7684
      11'd109  : in_data <= 14'h19da; // 'd6618
      11'd110  : in_data <= 14'h1caf; // 'd7343
      11'd111  : in_data <= 14'h0c67; // 'd3175
      11'd112  : in_data <= 14'h0cf5; // 'd3317
      11'd113  : in_data <= 14'h0249; // 'd585
      11'd114  : in_data <= 14'h089c; // 'd2204
      11'd115  : in_data <= 14'h151b; // 'd5403
      11'd116  : in_data <= 14'h021b; // 'd539
      11'd117  : in_data <= 14'h106a; // 'd4202
      11'd118  : in_data <= 14'h147e; // 'd5246
      11'd119  : in_data <= 14'h0315; // 'd789
      11'd120  : in_data <= 14'h0144; // 'd324
      11'd121  : in_data <= 14'h1bbd; // 'd7101
      11'd122  : in_data <= 14'h0b4f; // 'd2895
      11'd123  : in_data <= 14'h10f7; // 'd4343
      11'd124  : in_data <= 14'h0d30; // 'd3376
      11'd125  : in_data <= 14'h043f; // 'd1087
      11'd126  : in_data <= 14'h05b5; // 'd1461
      11'd127  : in_data <= 14'h0e92; // 'd3730
      11'd128  : in_data <= 14'h1c1a; // 'd7194
      11'd129  : in_data <= 14'h12b8; // 'd4792
      11'd130  : in_data <= 14'h0494; // 'd1172
      11'd131  : in_data <= 14'h161a; // 'd5658
      11'd132  : in_data <= 14'h104c; // 'd4172
      11'd133  : in_data <= 14'h0828; // 'd2088
      11'd134  : in_data <= 14'h095e; // 'd2398
      11'd135  : in_data <= 14'h1463; // 'd5219
      11'd136  : in_data <= 14'h1719; // 'd5913
      11'd137  : in_data <= 14'h0215; // 'd533
      11'd138  : in_data <= 14'h1a30; // 'd6704
      11'd139  : in_data <= 14'h0b95; // 'd2965
      11'd140  : in_data <= 14'h04e1; // 'd1249
      11'd141  : in_data <= 14'h0c10; // 'd3088
      11'd142  : in_data <= 14'h12bf; // 'd4799
      11'd143  : in_data <= 14'h15f2; // 'd5618
      11'd144  : in_data <= 14'h10c1; // 'd4289
      11'd145  : in_data <= 14'h05e1; // 'd1505
      11'd146  : in_data <= 14'h0cc2; // 'd3266
      11'd147  : in_data <= 14'h0f4f; // 'd3919
      11'd148  : in_data <= 14'h08ad; // 'd2221
      11'd149  : in_data <= 14'h151b; // 'd5403
      11'd150  : in_data <= 14'h005e; // 'd94
      11'd151  : in_data <= 14'h1a3e; // 'd6718
      11'd152  : in_data <= 14'h010e; // 'd270
      11'd153  : in_data <= 14'h1836; // 'd6198
      11'd154  : in_data <= 14'h18a6; // 'd6310
      11'd155  : in_data <= 14'h05eb; // 'd1515
      11'd156  : in_data <= 14'h1a40; // 'd6720
      11'd157  : in_data <= 14'h1267; // 'd4711
      11'd158  : in_data <= 14'h15cd; // 'd5581
      11'd159  : in_data <= 14'h145a; // 'd5210
      11'd160  : in_data <= 14'h073f; // 'd1855
      11'd161  : in_data <= 14'h1577; // 'd5495
      11'd162  : in_data <= 14'h1691; // 'd5777
      11'd163  : in_data <= 14'h0893; // 'd2195
      11'd164  : in_data <= 14'h087a; // 'd2170
      11'd165  : in_data <= 14'h0971; // 'd2417
      11'd166  : in_data <= 14'h114b; // 'd4427
      11'd167  : in_data <= 14'h1439; // 'd5177
      11'd168  : in_data <= 14'h10d0; // 'd4304
      11'd169  : in_data <= 14'h1bd3; // 'd7123
      11'd170  : in_data <= 14'h01ca; // 'd458
      11'd171  : in_data <= 14'h14a0; // 'd5280
      11'd172  : in_data <= 14'h1499; // 'd5273
      11'd173  : in_data <= 14'h15c1; // 'd5569
      11'd174  : in_data <= 14'h02a7; // 'd679
      11'd175  : in_data <= 14'h0900; // 'd2304
      11'd176  : in_data <= 14'h075a; // 'd1882
      11'd177  : in_data <= 14'h098e; // 'd2446
      11'd178  : in_data <= 14'h170b; // 'd5899
      11'd179  : in_data <= 14'h0867; // 'd2151
      11'd180  : in_data <= 14'h0f94; // 'd3988
      11'd181  : in_data <= 14'h0995; // 'd2453
      11'd182  : in_data <= 14'h1554; // 'd5460
      11'd183  : in_data <= 14'h0e7b; // 'd3707
      11'd184  : in_data <= 14'h02e0; // 'd736
      11'd185  : in_data <= 14'h1df2; // 'd7666
      11'd186  : in_data <= 14'h105b; // 'd4187
      11'd187  : in_data <= 14'h1a9e; // 'd6814
      11'd188  : in_data <= 14'h0910; // 'd2320
      11'd189  : in_data <= 14'h167b; // 'd5755
      11'd190  : in_data <= 14'h1dc7; // 'd7623
      11'd191  : in_data <= 14'h129b; // 'd4763
      11'd192  : in_data <= 14'h1aeb; // 'd6891
      11'd193  : in_data <= 14'h0d32; // 'd3378
      11'd194  : in_data <= 14'h1366; // 'd4966
      11'd195  : in_data <= 14'h19e9; // 'd6633
      11'd196  : in_data <= 14'h0719; // 'd1817
      11'd197  : in_data <= 14'h15c3; // 'd5571
      11'd198  : in_data <= 14'h122a; // 'd4650
      11'd199  : in_data <= 14'h03a4; // 'd932
      11'd200  : in_data <= 14'h01c5; // 'd453
      11'd201  : in_data <= 14'h0782; // 'd1922
      11'd202  : in_data <= 14'h13e8; // 'd5096
      11'd203  : in_data <= 14'h10b3; // 'd4275
      11'd204  : in_data <= 14'h08c8; // 'd2248
      11'd205  : in_data <= 14'h0fa7; // 'd4007
      11'd206  : in_data <= 14'h078e; // 'd1934
      11'd207  : in_data <= 14'h19a3; // 'd6563
      11'd208  : in_data <= 14'h04bf; // 'd1215
      11'd209  : in_data <= 14'h08f7; // 'd2295
      11'd210  : in_data <= 14'h1e59; // 'd7769
      11'd211  : in_data <= 14'h12e0; // 'd4832
      11'd212  : in_data <= 14'h0229; // 'd553
      11'd213  : in_data <= 14'h04c5; // 'd1221
      11'd214  : in_data <= 14'h11cc; // 'd4556
      11'd215  : in_data <= 14'h0321; // 'd801
      11'd216  : in_data <= 14'h0723; // 'd1827
      11'd217  : in_data <= 14'h03b0; // 'd944
      11'd218  : in_data <= 14'h160e; // 'd5646
      11'd219  : in_data <= 14'h1e1c; // 'd7708
      11'd220  : in_data <= 14'h0aca; // 'd2762
      11'd221  : in_data <= 14'h12e5; // 'd4837
      11'd222  : in_data <= 14'h032c; // 'd812
      11'd223  : in_data <= 14'h1104; // 'd4356
      11'd224  : in_data <= 14'h01ef; // 'd495
      11'd225  : in_data <= 14'h0fa0; // 'd4000
      11'd226  : in_data <= 14'h0f31; // 'd3889
      11'd227  : in_data <= 14'h189c; // 'd6300
      11'd228  : in_data <= 14'h0779; // 'd1913
      11'd229  : in_data <= 14'h11b7; // 'd4535
      11'd230  : in_data <= 14'h1e47; // 'd7751
      11'd231  : in_data <= 14'h00ac; // 'd172
      11'd232  : in_data <= 14'h15fe; // 'd5630
      11'd233  : in_data <= 14'h1515; // 'd5397
      11'd234  : in_data <= 14'h01cd; // 'd461
      11'd235  : in_data <= 14'h0af0; // 'd2800
      11'd236  : in_data <= 14'h0755; // 'd1877
      11'd237  : in_data <= 14'h087a; // 'd2170
      11'd238  : in_data <= 14'h02b2; // 'd690
      11'd239  : in_data <= 14'h0128; // 'd296
      11'd240  : in_data <= 14'h0c30; // 'd3120
      11'd241  : in_data <= 14'h1c61; // 'd7265
      11'd242  : in_data <= 14'h070c; // 'd1804
      11'd243  : in_data <= 14'h0d7e; // 'd3454
      11'd244  : in_data <= 14'h14f1; // 'd5361
      11'd245  : in_data <= 14'h0a51; // 'd2641
      11'd246  : in_data <= 14'h1940; // 'd6464
      11'd247  : in_data <= 14'h0b1e; // 'd2846
      11'd248  : in_data <= 14'h1d82; // 'd7554
      11'd249  : in_data <= 14'h0632; // 'd1586
      11'd250  : in_data <= 14'h17f6; // 'd6134
      11'd251  : in_data <= 14'h04b7; // 'd1207
      11'd252  : in_data <= 14'h1228; // 'd4648
      11'd253  : in_data <= 14'h0e45; // 'd3653
      11'd254  : in_data <= 14'h0abd; // 'd2749
      11'd255  : in_data <= 14'h0fdb; // 'd4059
      11'd256  : in_data <= 14'h1823; // 'd6179
      11'd257  : in_data <= 14'h18e4; // 'd6372
      11'd258  : in_data <= 14'h1374; // 'd4980
      11'd259  : in_data <= 14'h0d83; // 'd3459
      11'd260  : in_data <= 14'h0e0b; // 'd3595
      11'd261  : in_data <= 14'h1428; // 'd5160
      11'd262  : in_data <= 14'h0afc; // 'd2812
      11'd263  : in_data <= 14'h193c; // 'd6460
      11'd264  : in_data <= 14'h1ca6; // 'd7334
      11'd265  : in_data <= 14'h18d7; // 'd6359
      11'd266  : in_data <= 14'h1295; // 'd4757
      11'd267  : in_data <= 14'h1130; // 'd4400
      11'd268  : in_data <= 14'h0799; // 'd1945
      11'd269  : in_data <= 14'h1cec; // 'd7404
      11'd270  : in_data <= 14'h1c4e; // 'd7246
      11'd271  : in_data <= 14'h11a4; // 'd4516
      11'd272  : in_data <= 14'h12db; // 'd4827
      11'd273  : in_data <= 14'h162d; // 'd5677
      11'd274  : in_data <= 14'h065d; // 'd1629
      11'd275  : in_data <= 14'h153b; // 'd5435
      11'd276  : in_data <= 14'h147a; // 'd5242
      11'd277  : in_data <= 14'h14fb; // 'd5371
      11'd278  : in_data <= 14'h0915; // 'd2325
      11'd279  : in_data <= 14'h1982; // 'd6530
      11'd280  : in_data <= 14'h158e; // 'd5518
      11'd281  : in_data <= 14'h1e19; // 'd7705
      11'd282  : in_data <= 14'h0f29; // 'd3881
      11'd283  : in_data <= 14'h0b90; // 'd2960
      11'd284  : in_data <= 14'h15a6; // 'd5542
      11'd285  : in_data <= 14'h0d89; // 'd3465
      11'd286  : in_data <= 14'h095e; // 'd2398
      11'd287  : in_data <= 14'h1e52; // 'd7762
      11'd288  : in_data <= 14'h17f9; // 'd6137
      11'd289  : in_data <= 14'h0efe; // 'd3838
      11'd290  : in_data <= 14'h17cc; // 'd6092
      11'd291  : in_data <= 14'h0c78; // 'd3192
      11'd292  : in_data <= 14'h0547; // 'd1351
      11'd293  : in_data <= 14'h0d32; // 'd3378
      11'd294  : in_data <= 14'h09db; // 'd2523
      11'd295  : in_data <= 14'h1bb4; // 'd7092
      11'd296  : in_data <= 14'h169d; // 'd5789
      11'd297  : in_data <= 14'h17af; // 'd6063
      11'd298  : in_data <= 14'h16e4; // 'd5860
      11'd299  : in_data <= 14'h103d; // 'd4157
      11'd300  : in_data <= 14'h0126; // 'd294
      11'd301  : in_data <= 14'h11e1; // 'd4577
      11'd302  : in_data <= 14'h03d9; // 'd985
      11'd303  : in_data <= 14'h0c8e; // 'd3214
      11'd304  : in_data <= 14'h0f6d; // 'd3949
      11'd305  : in_data <= 14'h044c; // 'd1100
      11'd306  : in_data <= 14'h1ad9; // 'd6873
      11'd307  : in_data <= 14'h18c2; // 'd6338
      11'd308  : in_data <= 14'h09fd; // 'd2557
      11'd309  : in_data <= 14'h0bae; // 'd2990
      11'd310  : in_data <= 14'h0be2; // 'd3042
      11'd311  : in_data <= 14'h178d; // 'd6029
      11'd312  : in_data <= 14'h0e3b; // 'd3643
      11'd313  : in_data <= 14'h0adc; // 'd2780
      11'd314  : in_data <= 14'h01f5; // 'd501
      11'd315  : in_data <= 14'h0043; // 'd67
      11'd316  : in_data <= 14'h0919; // 'd2329
      11'd317  : in_data <= 14'h0c13; // 'd3091
      11'd318  : in_data <= 14'h0a8f; // 'd2703
      11'd319  : in_data <= 14'h13d5; // 'd5077
      11'd320  : in_data <= 14'h0e72; // 'd3698
      11'd321  : in_data <= 14'h122f; // 'd4655
      11'd322  : in_data <= 14'h0321; // 'd801
      11'd323  : in_data <= 14'h1b0f; // 'd6927
      11'd324  : in_data <= 14'h0548; // 'd1352
      11'd325  : in_data <= 14'h153f; // 'd5439
      11'd326  : in_data <= 14'h05d2; // 'd1490
      11'd327  : in_data <= 14'h0016; // 'd22
      11'd328  : in_data <= 14'h0f78; // 'd3960
      11'd329  : in_data <= 14'h1e4c; // 'd7756
      11'd330  : in_data <= 14'h1a4d; // 'd6733
      11'd331  : in_data <= 14'h1219; // 'd4633
      11'd332  : in_data <= 14'h175b; // 'd5979
      11'd333  : in_data <= 14'h0f3b; // 'd3899
      11'd334  : in_data <= 14'h10c6; // 'd4294
      11'd335  : in_data <= 14'h1adb; // 'd6875
      11'd336  : in_data <= 14'h13ae; // 'd5038
      11'd337  : in_data <= 14'h10e8; // 'd4328
      11'd338  : in_data <= 14'h0e69; // 'd3689
      11'd339  : in_data <= 14'h149d; // 'd5277
      11'd340  : in_data <= 14'h1573; // 'd5491
      11'd341  : in_data <= 14'h16aa; // 'd5802
      11'd342  : in_data <= 14'h0f3e; // 'd3902
      11'd343  : in_data <= 14'h081e; // 'd2078
      11'd344  : in_data <= 14'h1ac1; // 'd6849
      11'd345  : in_data <= 14'h0a4d; // 'd2637
      11'd346  : in_data <= 14'h01f0; // 'd496
      11'd347  : in_data <= 14'h0356; // 'd854
      11'd348  : in_data <= 14'h055a; // 'd1370
      11'd349  : in_data <= 14'h1c62; // 'd7266
      11'd350  : in_data <= 14'h0733; // 'd1843
      11'd351  : in_data <= 14'h1dc4; // 'd7620
      11'd352  : in_data <= 14'h08d7; // 'd2263
      11'd353  : in_data <= 14'h11c9; // 'd4553
      11'd354  : in_data <= 14'h1413; // 'd5139
      11'd355  : in_data <= 14'h0414; // 'd1044
      11'd356  : in_data <= 14'h11a5; // 'd4517
      11'd357  : in_data <= 14'h17a5; // 'd6053
      11'd358  : in_data <= 14'h10d6; // 'd4310
      11'd359  : in_data <= 14'h06fa; // 'd1786
      11'd360  : in_data <= 14'h0eee; // 'd3822
      11'd361  : in_data <= 14'h06b0; // 'd1712
      11'd362  : in_data <= 14'h1762; // 'd5986
      11'd363  : in_data <= 14'h0b0b; // 'd2827
      11'd364  : in_data <= 14'h022b; // 'd555
      11'd365  : in_data <= 14'h1238; // 'd4664
      11'd366  : in_data <= 14'h1bd4; // 'd7124
      11'd367  : in_data <= 14'h018c; // 'd396
      11'd368  : in_data <= 14'h0668; // 'd1640
      11'd369  : in_data <= 14'h12ad; // 'd4781
      11'd370  : in_data <= 14'h0c03; // 'd3075
      11'd371  : in_data <= 14'h17df; // 'd6111
      11'd372  : in_data <= 14'h1b52; // 'd6994
      11'd373  : in_data <= 14'h0bed; // 'd3053
      11'd374  : in_data <= 14'h1e49; // 'd7753
      11'd375  : in_data <= 14'h14d6; // 'd5334
      11'd376  : in_data <= 14'h0848; // 'd2120
      11'd377  : in_data <= 14'h0a1b; // 'd2587
      11'd378  : in_data <= 14'h190e; // 'd6414
      11'd379  : in_data <= 14'h0623; // 'd1571
      11'd380  : in_data <= 14'h1e43; // 'd7747
      11'd381  : in_data <= 14'h1c55; // 'd7253
      11'd382  : in_data <= 14'h1126; // 'd4390
      11'd383  : in_data <= 14'h122c; // 'd4652
      11'd384  : in_data <= 14'h18ab; // 'd6315
      11'd385  : in_data <= 14'h0b17; // 'd2839
      11'd386  : in_data <= 14'h1b24; // 'd6948
      11'd387  : in_data <= 14'h1e38; // 'd7736
      11'd388  : in_data <= 14'h168c; // 'd5772
      11'd389  : in_data <= 14'h0a6f; // 'd2671
      11'd390  : in_data <= 14'h156d; // 'd5485
      11'd391  : in_data <= 14'h1126; // 'd4390
      11'd392  : in_data <= 14'h0913; // 'd2323
      11'd393  : in_data <= 14'h17ff; // 'd6143
      11'd394  : in_data <= 14'h14a3; // 'd5283
      11'd395  : in_data <= 14'h0ae9; // 'd2793
      11'd396  : in_data <= 14'h19b0; // 'd6576
      11'd397  : in_data <= 14'h1023; // 'd4131
      11'd398  : in_data <= 14'h140f; // 'd5135
      11'd399  : in_data <= 14'h1e4e; // 'd7758
      11'd400  : in_data <= 14'h14c5; // 'd5317
      11'd401  : in_data <= 14'h1041; // 'd4161
      11'd402  : in_data <= 14'h0732; // 'd1842
      11'd403  : in_data <= 14'h17e3; // 'd6115
      11'd404  : in_data <= 14'h11ba; // 'd4538
      11'd405  : in_data <= 14'h121b; // 'd4635
      11'd406  : in_data <= 14'h0bb4; // 'd2996
      11'd407  : in_data <= 14'h07e1; // 'd2017
      11'd408  : in_data <= 14'h09b4; // 'd2484
      11'd409  : in_data <= 14'h1b22; // 'd6946
      11'd410  : in_data <= 14'h0a17; // 'd2583
      11'd411  : in_data <= 14'h0d84; // 'd3460
      11'd412  : in_data <= 14'h1992; // 'd6546
      11'd413  : in_data <= 14'h1002; // 'd4098
      11'd414  : in_data <= 14'h1b77; // 'd7031
      11'd415  : in_data <= 14'h0036; // 'd54
      11'd416  : in_data <= 14'h085b; // 'd2139
      11'd417  : in_data <= 14'h0d96; // 'd3478
      11'd418  : in_data <= 14'h0b7d; // 'd2941
      11'd419  : in_data <= 14'h161d; // 'd5661
      11'd420  : in_data <= 14'h0ec4; // 'd3780
      11'd421  : in_data <= 14'h0991; // 'd2449
      11'd422  : in_data <= 14'h0711; // 'd1809
      11'd423  : in_data <= 14'h020e; // 'd526
      11'd424  : in_data <= 14'h0a7d; // 'd2685
      11'd425  : in_data <= 14'h011b; // 'd283
      11'd426  : in_data <= 14'h0776; // 'd1910
      11'd427  : in_data <= 14'h0889; // 'd2185
      11'd428  : in_data <= 14'h140d; // 'd5133
      11'd429  : in_data <= 14'h1819; // 'd6169
      11'd430  : in_data <= 14'h1980; // 'd6528
      11'd431  : in_data <= 14'h102f; // 'd4143
      11'd432  : in_data <= 14'h06d8; // 'd1752
      11'd433  : in_data <= 14'h0868; // 'd2152
      11'd434  : in_data <= 14'h186e; // 'd6254
      11'd435  : in_data <= 14'h1c46; // 'd7238
      11'd436  : in_data <= 14'h1700; // 'd5888
      11'd437  : in_data <= 14'h1098; // 'd4248
      11'd438  : in_data <= 14'h1081; // 'd4225
      11'd439  : in_data <= 14'h0c30; // 'd3120
      11'd440  : in_data <= 14'h16a9; // 'd5801
      11'd441  : in_data <= 14'h0d50; // 'd3408
      11'd442  : in_data <= 14'h1148; // 'd4424
      11'd443  : in_data <= 14'h0c15; // 'd3093
      11'd444  : in_data <= 14'h0142; // 'd322
      11'd445  : in_data <= 14'h0fd1; // 'd4049
      11'd446  : in_data <= 14'h13b1; // 'd5041
      11'd447  : in_data <= 14'h1259; // 'd4697
      11'd448  : in_data <= 14'h114c; // 'd4428
      11'd449  : in_data <= 14'h1958; // 'd6488
      11'd450  : in_data <= 14'h034f; // 'd847
      11'd451  : in_data <= 14'h0eae; // 'd3758
      11'd452  : in_data <= 14'h109b; // 'd4251
      11'd453  : in_data <= 14'h1b33; // 'd6963
      11'd454  : in_data <= 14'h1147; // 'd4423
      11'd455  : in_data <= 14'h0b06; // 'd2822
      11'd456  : in_data <= 14'h11bb; // 'd4539
      11'd457  : in_data <= 14'h0d49; // 'd3401
      11'd458  : in_data <= 14'h16c2; // 'd5826
      11'd459  : in_data <= 14'h079f; // 'd1951
      11'd460  : in_data <= 14'h07b9; // 'd1977
      11'd461  : in_data <= 14'h1b29; // 'd6953
      11'd462  : in_data <= 14'h030a; // 'd778
      11'd463  : in_data <= 14'h11c3; // 'd4547
      11'd464  : in_data <= 14'h0bd2; // 'd3026
      11'd465  : in_data <= 14'h1124; // 'd4388
      11'd466  : in_data <= 14'h0569; // 'd1385
      11'd467  : in_data <= 14'h139c; // 'd5020
      11'd468  : in_data <= 14'h09d3; // 'd2515
      11'd469  : in_data <= 14'h19c3; // 'd6595
      11'd470  : in_data <= 14'h14a4; // 'd5284
      11'd471  : in_data <= 14'h11dd; // 'd4573
      11'd472  : in_data <= 14'h0a81; // 'd2689
      11'd473  : in_data <= 14'h165d; // 'd5725
      11'd474  : in_data <= 14'h1715; // 'd5909
      11'd475  : in_data <= 14'h1121; // 'd4385
      11'd476  : in_data <= 14'h0777; // 'd1911
      11'd477  : in_data <= 14'h09bb; // 'd2491
      11'd478  : in_data <= 14'h1a6c; // 'd6764
      11'd479  : in_data <= 14'h0297; // 'd663
      11'd480  : in_data <= 14'h0682; // 'd1666
      11'd481  : in_data <= 14'h0d7e; // 'd3454
      11'd482  : in_data <= 14'h0a6a; // 'd2666
      11'd483  : in_data <= 14'h04b0; // 'd1200
      11'd484  : in_data <= 14'h176e; // 'd5998
      11'd485  : in_data <= 14'h18e3; // 'd6371
      11'd486  : in_data <= 14'h0b79; // 'd2937
      11'd487  : in_data <= 14'h173d; // 'd5949
      11'd488  : in_data <= 14'h115d; // 'd4445
      11'd489  : in_data <= 14'h0ecd; // 'd3789
      11'd490  : in_data <= 14'h1d9f; // 'd7583
      11'd491  : in_data <= 14'h104e; // 'd4174
      11'd492  : in_data <= 14'h0442; // 'd1090
      11'd493  : in_data <= 14'h07f7; // 'd2039
      11'd494  : in_data <= 14'h08be; // 'd2238
      11'd495  : in_data <= 14'h0e55; // 'd3669
      11'd496  : in_data <= 14'h1350; // 'd4944
      11'd497  : in_data <= 14'h0b0a; // 'd2826
      11'd498  : in_data <= 14'h02ba; // 'd698
      11'd499  : in_data <= 14'h14a8; // 'd5288
      11'd500  : in_data <= 14'h047a; // 'd1146
      11'd501  : in_data <= 14'h1da0; // 'd7584
      11'd502  : in_data <= 14'h062c; // 'd1580
      11'd503  : in_data <= 14'h1369; // 'd4969
      11'd504  : in_data <= 14'h06bb; // 'd1723
      11'd505  : in_data <= 14'h1cb2; // 'd7346
      11'd506  : in_data <= 14'h18a9; // 'd6313
      11'd507  : in_data <= 14'h1b65; // 'd7013
      11'd508  : in_data <= 14'h07b0; // 'd1968
      11'd509  : in_data <= 14'h0d51; // 'd3409
      11'd510  : in_data <= 14'h11e9; // 'd4585
      11'd511  : in_data <= 14'h18a3; // 'd6307
      11'd512  : in_data <= 14'h1e19; // 'd7705
      11'd513  : in_data <= 14'h1a63; // 'd6755
      11'd514  : in_data <= 14'h1a31; // 'd6705
      11'd515  : in_data <= 14'h12ca; // 'd4810
      11'd516  : in_data <= 14'h0061; // 'd97
      11'd517  : in_data <= 14'h0647; // 'd1607
      11'd518  : in_data <= 14'h0a40; // 'd2624
      11'd519  : in_data <= 14'h1b75; // 'd7029
      11'd520  : in_data <= 14'h02df; // 'd735
      11'd521  : in_data <= 14'h1c35; // 'd7221
      11'd522  : in_data <= 14'h04a4; // 'd1188
      11'd523  : in_data <= 14'h0115; // 'd277
      11'd524  : in_data <= 14'h0457; // 'd1111
      11'd525  : in_data <= 14'h02f0; // 'd752
      11'd526  : in_data <= 14'h0984; // 'd2436
      11'd527  : in_data <= 14'h0d74; // 'd3444
      11'd528  : in_data <= 14'h16c3; // 'd5827
      11'd529  : in_data <= 14'h0875; // 'd2165
      11'd530  : in_data <= 14'h19d2; // 'd6610
      11'd531  : in_data <= 14'h0de3; // 'd3555
      11'd532  : in_data <= 14'h08a0; // 'd2208
      11'd533  : in_data <= 14'h19f2; // 'd6642
      11'd534  : in_data <= 14'h008a; // 'd138
      11'd535  : in_data <= 14'h10fc; // 'd4348
      11'd536  : in_data <= 14'h0850; // 'd2128
      11'd537  : in_data <= 14'h0885; // 'd2181
      11'd538  : in_data <= 14'h1583; // 'd5507
      11'd539  : in_data <= 14'h0db5; // 'd3509
      11'd540  : in_data <= 14'h1358; // 'd4952
      11'd541  : in_data <= 14'h0c4b; // 'd3147
      11'd542  : in_data <= 14'h121b; // 'd4635
      11'd543  : in_data <= 14'h12bd; // 'd4797
      11'd544  : in_data <= 14'h1d28; // 'd7464
      11'd545  : in_data <= 14'h0eb6; // 'd3766
      11'd546  : in_data <= 14'h0337; // 'd823
      11'd547  : in_data <= 14'h00f3; // 'd243
      11'd548  : in_data <= 14'h0aeb; // 'd2795
      11'd549  : in_data <= 14'h0569; // 'd1385
      11'd550  : in_data <= 14'h0e91; // 'd3729
      11'd551  : in_data <= 14'h0a9d; // 'd2717
      11'd552  : in_data <= 14'h05ef; // 'd1519
      11'd553  : in_data <= 14'h1965; // 'd6501
      11'd554  : in_data <= 14'h0aab; // 'd2731
      11'd555  : in_data <= 14'h1481; // 'd5249
      11'd556  : in_data <= 14'h0132; // 'd306
      11'd557  : in_data <= 14'h019d; // 'd413
      11'd558  : in_data <= 14'h17cd; // 'd6093
      11'd559  : in_data <= 14'h1e66; // 'd7782
      11'd560  : in_data <= 14'h0bb9; // 'd3001
      11'd561  : in_data <= 14'h15d5; // 'd5589
      11'd562  : in_data <= 14'h1d3e; // 'd7486
      11'd563  : in_data <= 14'h0b78; // 'd2936
      11'd564  : in_data <= 14'h0f93; // 'd3987
      11'd565  : in_data <= 14'h1e4d; // 'd7757
      11'd566  : in_data <= 14'h12a5; // 'd4773
      11'd567  : in_data <= 14'h1a1e; // 'd6686
      11'd568  : in_data <= 14'h090c; // 'd2316
      11'd569  : in_data <= 14'h1e83; // 'd7811
      11'd570  : in_data <= 14'h11fd; // 'd4605
      11'd571  : in_data <= 14'h08e1; // 'd2273
      11'd572  : in_data <= 14'h0802; // 'd2050
      11'd573  : in_data <= 14'h0ad9; // 'd2777
      11'd574  : in_data <= 14'h0c2c; // 'd3116
      11'd575  : in_data <= 14'h17f3; // 'd6131
      11'd576  : in_data <= 14'h0a8c; // 'd2700
      11'd577  : in_data <= 14'h10f3; // 'd4339
      11'd578  : in_data <= 14'h010c; // 'd268
      11'd579  : in_data <= 14'h05c3; // 'd1475
      11'd580  : in_data <= 14'h04f4; // 'd1268
      11'd581  : in_data <= 14'h04b0; // 'd1200
      11'd582  : in_data <= 14'h160a; // 'd5642
      11'd583  : in_data <= 14'h1e1f; // 'd7711
      11'd584  : in_data <= 14'h1b9a; // 'd7066
      11'd585  : in_data <= 14'h1d0f; // 'd7439
      11'd586  : in_data <= 14'h09c1; // 'd2497
      11'd587  : in_data <= 14'h0374; // 'd884
      11'd588  : in_data <= 14'h1774; // 'd6004
      11'd589  : in_data <= 14'h1cac; // 'd7340
      11'd590  : in_data <= 14'h1230; // 'd4656
      11'd591  : in_data <= 14'h02a2; // 'd674
      11'd592  : in_data <= 14'h01c8; // 'd456
      11'd593  : in_data <= 14'h1713; // 'd5907
      11'd594  : in_data <= 14'h0a07; // 'd2567
      11'd595  : in_data <= 14'h0449; // 'd1097
      11'd596  : in_data <= 14'h0d0e; // 'd3342
      11'd597  : in_data <= 14'h0aa8; // 'd2728
      11'd598  : in_data <= 14'h17a8; // 'd6056
      11'd599  : in_data <= 14'h0000; // 'd0
      11'd600  : in_data <= 14'h0477; // 'd1143
      11'd601  : in_data <= 14'h0046; // 'd70
      11'd602  : in_data <= 14'h0221; // 'd545
      11'd603  : in_data <= 14'h1bc7; // 'd7111
      11'd604  : in_data <= 14'h0069; // 'd105
      11'd605  : in_data <= 14'h1b0f; // 'd6927
      11'd606  : in_data <= 14'h1d5e; // 'd7518
      11'd607  : in_data <= 14'h06af; // 'd1711
      11'd608  : in_data <= 14'h0940; // 'd2368
      11'd609  : in_data <= 14'h0b47; // 'd2887
      11'd610  : in_data <= 14'h1ce4; // 'd7396
      11'd611  : in_data <= 14'h036c; // 'd876
      11'd612  : in_data <= 14'h0263; // 'd611
      11'd613  : in_data <= 14'h115a; // 'd4442
      11'd614  : in_data <= 14'h13e1; // 'd5089
      11'd615  : in_data <= 14'h176f; // 'd5999
      11'd616  : in_data <= 14'h05de; // 'd1502
      11'd617  : in_data <= 14'h0ac8; // 'd2760
      11'd618  : in_data <= 14'h1af2; // 'd6898
      11'd619  : in_data <= 14'h0492; // 'd1170
      11'd620  : in_data <= 14'h0804; // 'd2052
      11'd621  : in_data <= 14'h1078; // 'd4216
      11'd622  : in_data <= 14'h10af; // 'd4271
      11'd623  : in_data <= 14'h0209; // 'd521
      11'd624  : in_data <= 14'h17eb; // 'd6123
      11'd625  : in_data <= 14'h0af9; // 'd2809
      11'd626  : in_data <= 14'h0b7f; // 'd2943
      11'd627  : in_data <= 14'h09d6; // 'd2518
      11'd628  : in_data <= 14'h04d7; // 'd1239
      11'd629  : in_data <= 14'h008e; // 'd142
      11'd630  : in_data <= 14'h158e; // 'd5518
      11'd631  : in_data <= 14'h1b7a; // 'd7034
      11'd632  : in_data <= 14'h1b69; // 'd7017
      11'd633  : in_data <= 14'h146c; // 'd5228
      11'd634  : in_data <= 14'h00ec; // 'd236
      11'd635  : in_data <= 14'h0a80; // 'd2688
      11'd636  : in_data <= 14'h0e66; // 'd3686
      11'd637  : in_data <= 14'h1057; // 'd4183
      11'd638  : in_data <= 14'h018e; // 'd398
      11'd639  : in_data <= 14'h05b7; // 'd1463
      11'd640  : in_data <= 14'h0538; // 'd1336
      11'd641  : in_data <= 14'h080c; // 'd2060
      11'd642  : in_data <= 14'h0f5e; // 'd3934
      11'd643  : in_data <= 14'h120a; // 'd4618
      11'd644  : in_data <= 14'h04bb; // 'd1211
      11'd645  : in_data <= 14'h18f0; // 'd6384
      11'd646  : in_data <= 14'h0de1; // 'd3553
      11'd647  : in_data <= 14'h11ca; // 'd4554
      11'd648  : in_data <= 14'h18d6; // 'd6358
      11'd649  : in_data <= 14'h100e; // 'd4110
      11'd650  : in_data <= 14'h1878; // 'd6264
      11'd651  : in_data <= 14'h0b2d; // 'd2861
      11'd652  : in_data <= 14'h1ad0; // 'd6864
      11'd653  : in_data <= 14'h1e7a; // 'd7802
      11'd654  : in_data <= 14'h0d5b; // 'd3419
      11'd655  : in_data <= 14'h14d1; // 'd5329
      11'd656  : in_data <= 14'h0d05; // 'd3333
      11'd657  : in_data <= 14'h0f25; // 'd3877
      11'd658  : in_data <= 14'h0d79; // 'd3449
      11'd659  : in_data <= 14'h1330; // 'd4912
      11'd660  : in_data <= 14'h0db7; // 'd3511
      11'd661  : in_data <= 14'h0ac4; // 'd2756
      11'd662  : in_data <= 14'h1035; // 'd4149
      11'd663  : in_data <= 14'h0f56; // 'd3926
      11'd664  : in_data <= 14'h1cdd; // 'd7389
      11'd665  : in_data <= 14'h0aa7; // 'd2727
      11'd666  : in_data <= 14'h1009; // 'd4105
      11'd667  : in_data <= 14'h0a7a; // 'd2682
      11'd668  : in_data <= 14'h0f6f; // 'd3951
      11'd669  : in_data <= 14'h17f8; // 'd6136
      11'd670  : in_data <= 14'h058d; // 'd1421
      11'd671  : in_data <= 14'h1d1c; // 'd7452
      11'd672  : in_data <= 14'h1607; // 'd5639
      11'd673  : in_data <= 14'h1b42; // 'd6978
      11'd674  : in_data <= 14'h12f3; // 'd4851
      11'd675  : in_data <= 14'h0b2e; // 'd2862
      11'd676  : in_data <= 14'h16f7; // 'd5879
      11'd677  : in_data <= 14'h1a3e; // 'd6718
      11'd678  : in_data <= 14'h03af; // 'd943
      11'd679  : in_data <= 14'h01c9; // 'd457
      11'd680  : in_data <= 14'h04fe; // 'd1278
      11'd681  : in_data <= 14'h018e; // 'd398
      11'd682  : in_data <= 14'h106b; // 'd4203
      11'd683  : in_data <= 14'h14a9; // 'd5289
      11'd684  : in_data <= 14'h0310; // 'd784
      11'd685  : in_data <= 14'h0974; // 'd2420
      11'd686  : in_data <= 14'h1295; // 'd4757
      11'd687  : in_data <= 14'h1144; // 'd4420
      11'd688  : in_data <= 14'h02cd; // 'd717
      11'd689  : in_data <= 14'h07a6; // 'd1958
      11'd690  : in_data <= 14'h0d1b; // 'd3355
      11'd691  : in_data <= 14'h019f; // 'd415
      11'd692  : in_data <= 14'h052c; // 'd1324
      11'd693  : in_data <= 14'h16b0; // 'd5808
      11'd694  : in_data <= 14'h111d; // 'd4381
      11'd695  : in_data <= 14'h06db; // 'd1755
      11'd696  : in_data <= 14'h035e; // 'd862
      11'd697  : in_data <= 14'h0d74; // 'd3444
      11'd698  : in_data <= 14'h0b16; // 'd2838
      11'd699  : in_data <= 14'h02c1; // 'd705
      11'd700  : in_data <= 14'h1aeb; // 'd6891
      11'd701  : in_data <= 14'h0cdc; // 'd3292
      11'd702  : in_data <= 14'h1e7c; // 'd7804
      11'd703  : in_data <= 14'h0d76; // 'd3446
      11'd704  : in_data <= 14'h07fa; // 'd2042
      11'd705  : in_data <= 14'h0adf; // 'd2783
      11'd706  : in_data <= 14'h1528; // 'd5416
      11'd707  : in_data <= 14'h0c4f; // 'd3151
      11'd708  : in_data <= 14'h162b; // 'd5675
      11'd709  : in_data <= 14'h17d9; // 'd6105
      11'd710  : in_data <= 14'h04e1; // 'd1249
      11'd711  : in_data <= 14'h0d7b; // 'd3451
      11'd712  : in_data <= 14'h1bc9; // 'd7113
      11'd713  : in_data <= 14'h1445; // 'd5189
      11'd714  : in_data <= 14'h1704; // 'd5892
      11'd715  : in_data <= 14'h1b40; // 'd6976
      11'd716  : in_data <= 14'h1613; // 'd5651
      11'd717  : in_data <= 14'h1e7b; // 'd7803
      11'd718  : in_data <= 14'h0e4e; // 'd3662
      11'd719  : in_data <= 14'h1a08; // 'd6664
      11'd720  : in_data <= 14'h1ce4; // 'd7396
      11'd721  : in_data <= 14'h0129; // 'd297
      11'd722  : in_data <= 14'h1abf; // 'd6847
      11'd723  : in_data <= 14'h1b99; // 'd7065
      11'd724  : in_data <= 14'h1c25; // 'd7205
      11'd725  : in_data <= 14'h051d; // 'd1309
      11'd726  : in_data <= 14'h1310; // 'd4880
      11'd727  : in_data <= 14'h0307; // 'd775
      11'd728  : in_data <= 14'h0ccd; // 'd3277
      11'd729  : in_data <= 14'h11be; // 'd4542
      11'd730  : in_data <= 14'h192e; // 'd6446
      11'd731  : in_data <= 14'h1012; // 'd4114
      11'd732  : in_data <= 14'h1e0a; // 'd7690
      11'd733  : in_data <= 14'h1693; // 'd5779
      11'd734  : in_data <= 14'h1502; // 'd5378
      11'd735  : in_data <= 14'h1943; // 'd6467
      11'd736  : in_data <= 14'h1689; // 'd5769
      11'd737  : in_data <= 14'h1958; // 'd6488
      11'd738  : in_data <= 14'h193d; // 'd6461
      11'd739  : in_data <= 14'h146d; // 'd5229
      11'd740  : in_data <= 14'h1bdc; // 'd7132
      11'd741  : in_data <= 14'h1723; // 'd5923
      11'd742  : in_data <= 14'h11b5; // 'd4533
      11'd743  : in_data <= 14'h12c5; // 'd4805
      11'd744  : in_data <= 14'h14ff; // 'd5375
      11'd745  : in_data <= 14'h1299; // 'd4761
      11'd746  : in_data <= 14'h0aa8; // 'd2728
      11'd747  : in_data <= 14'h17f4; // 'd6132
      11'd748  : in_data <= 14'h114d; // 'd4429
      11'd749  : in_data <= 14'h1bd0; // 'd7120
      11'd750  : in_data <= 14'h05d5; // 'd1493
      11'd751  : in_data <= 14'h1d40; // 'd7488
      11'd752  : in_data <= 14'h0a29; // 'd2601
      11'd753  : in_data <= 14'h01ab; // 'd427
      11'd754  : in_data <= 14'h0f88; // 'd3976
      11'd755  : in_data <= 14'h069e; // 'd1694
      11'd756  : in_data <= 14'h1b86; // 'd7046
      11'd757  : in_data <= 14'h17d4; // 'd6100
      11'd758  : in_data <= 14'h0265; // 'd613
      11'd759  : in_data <= 14'h0828; // 'd2088
      11'd760  : in_data <= 14'h016c; // 'd364
      11'd761  : in_data <= 14'h10ba; // 'd4282
      11'd762  : in_data <= 14'h1e5f; // 'd7775
      11'd763  : in_data <= 14'h0fe4; // 'd4068
      11'd764  : in_data <= 14'h121b; // 'd4635
      11'd765  : in_data <= 14'h0e47; // 'd3655
      11'd766  : in_data <= 14'h0d00; // 'd3328
      11'd767  : in_data <= 14'h172c; // 'd5932
      11'd768  : in_data <= 14'h0d6b; // 'd3435
      11'd769  : in_data <= 14'h0d31; // 'd3377
      11'd770  : in_data <= 14'h0816; // 'd2070
      11'd771  : in_data <= 14'h173e; // 'd5950
      11'd772  : in_data <= 14'h1da4; // 'd7588
      11'd773  : in_data <= 14'h0338; // 'd824
      11'd774  : in_data <= 14'h0889; // 'd2185
      11'd775  : in_data <= 14'h023e; // 'd574
      11'd776  : in_data <= 14'h081c; // 'd2076
      11'd777  : in_data <= 14'h0052; // 'd82
      11'd778  : in_data <= 14'h0c14; // 'd3092
      11'd779  : in_data <= 14'h0fd4; // 'd4052
      11'd780  : in_data <= 14'h1c1e; // 'd7198
      11'd781  : in_data <= 14'h1ba0; // 'd7072
      11'd782  : in_data <= 14'h1b28; // 'd6952
      11'd783  : in_data <= 14'h15c0; // 'd5568
      11'd784  : in_data <= 14'h1b0d; // 'd6925
      11'd785  : in_data <= 14'h02ca; // 'd714
      11'd786  : in_data <= 14'h043d; // 'd1085
      11'd787  : in_data <= 14'h02cc; // 'd716
      11'd788  : in_data <= 14'h12f1; // 'd4849
      11'd789  : in_data <= 14'h15bb; // 'd5563
      11'd790  : in_data <= 14'h1e62; // 'd7778
      11'd791  : in_data <= 14'h0dda; // 'd3546
      11'd792  : in_data <= 14'h07f4; // 'd2036
      11'd793  : in_data <= 14'h150b; // 'd5387
      11'd794  : in_data <= 14'h16ad; // 'd5805
      11'd795  : in_data <= 14'h17d2; // 'd6098
      11'd796  : in_data <= 14'h06e6; // 'd1766
      11'd797  : in_data <= 14'h0319; // 'd793
      11'd798  : in_data <= 14'h1278; // 'd4728
      11'd799  : in_data <= 14'h01ca; // 'd458
      11'd800  : in_data <= 14'h07ec; // 'd2028
      11'd801  : in_data <= 14'h1958; // 'd6488
      11'd802  : in_data <= 14'h13e3; // 'd5091
      11'd803  : in_data <= 14'h0603; // 'd1539
      11'd804  : in_data <= 14'h09ad; // 'd2477
      11'd805  : in_data <= 14'h19fa; // 'd6650
      11'd806  : in_data <= 14'h027d; // 'd637
      11'd807  : in_data <= 14'h08e2; // 'd2274
      11'd808  : in_data <= 14'h1042; // 'd4162
      11'd809  : in_data <= 14'h11c3; // 'd4547
      11'd810  : in_data <= 14'h0c1f; // 'd3103
      11'd811  : in_data <= 14'h12f9; // 'd4857
      11'd812  : in_data <= 14'h08c4; // 'd2244
      11'd813  : in_data <= 14'h14c7; // 'd5319
      11'd814  : in_data <= 14'h08e8; // 'd2280
      11'd815  : in_data <= 14'h17f4; // 'd6132
      11'd816  : in_data <= 14'h19a4; // 'd6564
      11'd817  : in_data <= 14'h1525; // 'd5413
      11'd818  : in_data <= 14'h13ce; // 'd5070
      11'd819  : in_data <= 14'h0d3a; // 'd3386
      11'd820  : in_data <= 14'h1af3; // 'd6899
      11'd821  : in_data <= 14'h0b51; // 'd2897
      11'd822  : in_data <= 14'h124e; // 'd4686
      11'd823  : in_data <= 14'h067a; // 'd1658
      11'd824  : in_data <= 14'h16a8; // 'd5800
      11'd825  : in_data <= 14'h149b; // 'd5275
      11'd826  : in_data <= 14'h0b40; // 'd2880
      11'd827  : in_data <= 14'h006a; // 'd106
      11'd828  : in_data <= 14'h0e37; // 'd3639
      11'd829  : in_data <= 14'h1eaa; // 'd7850
      11'd830  : in_data <= 14'h1d62; // 'd7522
      11'd831  : in_data <= 14'h01b0; // 'd432
      11'd832  : in_data <= 14'h077f; // 'd1919
      11'd833  : in_data <= 14'h1cb1; // 'd7345
      11'd834  : in_data <= 14'h0af9; // 'd2809
      11'd835  : in_data <= 14'h1371; // 'd4977
      11'd836  : in_data <= 14'h1887; // 'd6279
      11'd837  : in_data <= 14'h062d; // 'd1581
      11'd838  : in_data <= 14'h03d9; // 'd985
      11'd839  : in_data <= 14'h029a; // 'd666
      11'd840  : in_data <= 14'h0bab; // 'd2987
      11'd841  : in_data <= 14'h121c; // 'd4636
      11'd842  : in_data <= 14'h0641; // 'd1601
      11'd843  : in_data <= 14'h1932; // 'd6450
      11'd844  : in_data <= 14'h0656; // 'd1622
      11'd845  : in_data <= 14'h0b18; // 'd2840
      11'd846  : in_data <= 14'h0407; // 'd1031
      11'd847  : in_data <= 14'h05a2; // 'd1442
      11'd848  : in_data <= 14'h0aa8; // 'd2728
      11'd849  : in_data <= 14'h1823; // 'd6179
      11'd850  : in_data <= 14'h11f4; // 'd4596
      11'd851  : in_data <= 14'h01f5; // 'd501
      11'd852  : in_data <= 14'h194b; // 'd6475
      11'd853  : in_data <= 14'h0d92; // 'd3474
      11'd854  : in_data <= 14'h1804; // 'd6148
      11'd855  : in_data <= 14'h1939; // 'd6457
      11'd856  : in_data <= 14'h074d; // 'd1869
      11'd857  : in_data <= 14'h1774; // 'd6004
      11'd858  : in_data <= 14'h04a5; // 'd1189
      11'd859  : in_data <= 14'h19e3; // 'd6627
      11'd860  : in_data <= 14'h122c; // 'd4652
      11'd861  : in_data <= 14'h17b9; // 'd6073
      11'd862  : in_data <= 14'h0a57; // 'd2647
      11'd863  : in_data <= 14'h1c15; // 'd7189
      11'd864  : in_data <= 14'h08ff; // 'd2303
      11'd865  : in_data <= 14'h16f1; // 'd5873
      11'd866  : in_data <= 14'h060e; // 'd1550
      11'd867  : in_data <= 14'h0ffc; // 'd4092
      11'd868  : in_data <= 14'h1057; // 'd4183
      11'd869  : in_data <= 14'h165c; // 'd5724
      11'd870  : in_data <= 14'h0203; // 'd515
      11'd871  : in_data <= 14'h18b3; // 'd6323
      11'd872  : in_data <= 14'h018c; // 'd396
      11'd873  : in_data <= 14'h02b8; // 'd696
      11'd874  : in_data <= 14'h1c2f; // 'd7215
      11'd875  : in_data <= 14'h1cec; // 'd7404
      11'd876  : in_data <= 14'h1b36; // 'd6966
      11'd877  : in_data <= 14'h1405; // 'd5125
      11'd878  : in_data <= 14'h06a8; // 'd1704
      11'd879  : in_data <= 14'h1ea2; // 'd7842
      11'd880  : in_data <= 14'h145e; // 'd5214
      11'd881  : in_data <= 14'h1a79; // 'd6777
      11'd882  : in_data <= 14'h1568; // 'd5480
      11'd883  : in_data <= 14'h136c; // 'd4972
      11'd884  : in_data <= 14'h02de; // 'd734
      11'd885  : in_data <= 14'h1e89; // 'd7817
      11'd886  : in_data <= 14'h1642; // 'd5698
      11'd887  : in_data <= 14'h0a62; // 'd2658
      11'd888  : in_data <= 14'h0ac1; // 'd2753
      11'd889  : in_data <= 14'h0e81; // 'd3713
      11'd890  : in_data <= 14'h177f; // 'd6015
      11'd891  : in_data <= 14'h0de9; // 'd3561
      11'd892  : in_data <= 14'h077a; // 'd1914
      11'd893  : in_data <= 14'h0932; // 'd2354
      11'd894  : in_data <= 14'h1e0c; // 'd7692
      11'd895  : in_data <= 14'h17b0; // 'd6064
      11'd896  : in_data <= 14'h0157; // 'd343
      11'd897  : in_data <= 14'h0e06; // 'd3590
      11'd898  : in_data <= 14'h057b; // 'd1403
      11'd899  : in_data <= 14'h113d; // 'd4413
      11'd900  : in_data <= 14'h081e; // 'd2078
      11'd901  : in_data <= 14'h1491; // 'd5265
      11'd902  : in_data <= 14'h08fc; // 'd2300
      11'd903  : in_data <= 14'h0fc6; // 'd4038
      11'd904  : in_data <= 14'h0e93; // 'd3731
      11'd905  : in_data <= 14'h182e; // 'd6190
      11'd906  : in_data <= 14'h1498; // 'd5272
      11'd907  : in_data <= 14'h1e0b; // 'd7691
      11'd908  : in_data <= 14'h1c78; // 'd7288
      11'd909  : in_data <= 14'h1b87; // 'd7047
      11'd910  : in_data <= 14'h1dce; // 'd7630
      11'd911  : in_data <= 14'h1465; // 'd5221
      11'd912  : in_data <= 14'h101c; // 'd4124
      11'd913  : in_data <= 14'h1169; // 'd4457
      11'd914  : in_data <= 14'h0886; // 'd2182
      11'd915  : in_data <= 14'h1c03; // 'd7171
      11'd916  : in_data <= 14'h0d49; // 'd3401
      11'd917  : in_data <= 14'h1da6; // 'd7590
      11'd918  : in_data <= 14'h03eb; // 'd1003
      11'd919  : in_data <= 14'h076f; // 'd1903
      11'd920  : in_data <= 14'h104c; // 'd4172
      11'd921  : in_data <= 14'h0864; // 'd2148
      11'd922  : in_data <= 14'h0176; // 'd374
      11'd923  : in_data <= 14'h01dd; // 'd477
      11'd924  : in_data <= 14'h0203; // 'd515
      11'd925  : in_data <= 14'h1407; // 'd5127
      11'd926  : in_data <= 14'h1ae4; // 'd6884
      11'd927  : in_data <= 14'h1562; // 'd5474
      11'd928  : in_data <= 14'h0af3; // 'd2803
      11'd929  : in_data <= 14'h0743; // 'd1859
      11'd930  : in_data <= 14'h15e6; // 'd5606
      11'd931  : in_data <= 14'h1d86; // 'd7558
      11'd932  : in_data <= 14'h05bd; // 'd1469
      11'd933  : in_data <= 14'h0ea5; // 'd3749
      11'd934  : in_data <= 14'h0178; // 'd376
      11'd935  : in_data <= 14'h124d; // 'd4685
      11'd936  : in_data <= 14'h1caf; // 'd7343
      11'd937  : in_data <= 14'h081d; // 'd2077
      11'd938  : in_data <= 14'h0299; // 'd665
      11'd939  : in_data <= 14'h0d1d; // 'd3357
      11'd940  : in_data <= 14'h00d4; // 'd212
      11'd941  : in_data <= 14'h0471; // 'd1137
      11'd942  : in_data <= 14'h016e; // 'd366
      11'd943  : in_data <= 14'h175b; // 'd5979
      11'd944  : in_data <= 14'h0931; // 'd2353
      11'd945  : in_data <= 14'h1758; // 'd5976
      11'd946  : in_data <= 14'h0861; // 'd2145
      11'd947  : in_data <= 14'h04d9; // 'd1241
      11'd948  : in_data <= 14'h15ae; // 'd5550
      11'd949  : in_data <= 14'h01e4; // 'd484
      11'd950  : in_data <= 14'h19c2; // 'd6594
      11'd951  : in_data <= 14'h03a7; // 'd935
      11'd952  : in_data <= 14'h13e1; // 'd5089
      11'd953  : in_data <= 14'h1ab3; // 'd6835
      11'd954  : in_data <= 14'h100b; // 'd4107
      11'd955  : in_data <= 14'h0abb; // 'd2747
      11'd956  : in_data <= 14'h0a57; // 'd2647
      11'd957  : in_data <= 14'h1e6c; // 'd7788
      11'd958  : in_data <= 14'h18ca; // 'd6346
      11'd959  : in_data <= 14'h0cd6; // 'd3286
      11'd960  : in_data <= 14'h0459; // 'd1113
      11'd961  : in_data <= 14'h01da; // 'd474
      11'd962  : in_data <= 14'h06e1; // 'd1761
      11'd963  : in_data <= 14'h0e91; // 'd3729
      11'd964  : in_data <= 14'h17d0; // 'd6096
      11'd965  : in_data <= 14'h014d; // 'd333
      11'd966  : in_data <= 14'h1c96; // 'd7318
      11'd967  : in_data <= 14'h063f; // 'd1599
      11'd968  : in_data <= 14'h0aea; // 'd2794
      11'd969  : in_data <= 14'h0748; // 'd1864
      11'd970  : in_data <= 14'h01a8; // 'd424
      11'd971  : in_data <= 14'h1a30; // 'd6704
      11'd972  : in_data <= 14'h181c; // 'd6172
      11'd973  : in_data <= 14'h06ea; // 'd1770
      11'd974  : in_data <= 14'h138d; // 'd5005
      11'd975  : in_data <= 14'h182f; // 'd6191
      11'd976  : in_data <= 14'h0ef0; // 'd3824
      11'd977  : in_data <= 14'h1183; // 'd4483
      11'd978  : in_data <= 14'h124b; // 'd4683
      11'd979  : in_data <= 14'h14f1; // 'd5361
      11'd980  : in_data <= 14'h15e1; // 'd5601
      11'd981  : in_data <= 14'h0e27; // 'd3623
      11'd982  : in_data <= 14'h080e; // 'd2062
      11'd983  : in_data <= 14'h0a2c; // 'd2604
      11'd984  : in_data <= 14'h1ec4; // 'd7876
      11'd985  : in_data <= 14'h0ef4; // 'd3828
      11'd986  : in_data <= 14'h1d21; // 'd7457
      11'd987  : in_data <= 14'h1978; // 'd6520
      11'd988  : in_data <= 14'h039f; // 'd927
      11'd989  : in_data <= 14'h0246; // 'd582
      11'd990  : in_data <= 14'h183c; // 'd6204
      11'd991  : in_data <= 14'h13e3; // 'd5091
      11'd992  : in_data <= 14'h1333; // 'd4915
      11'd993  : in_data <= 14'h0677; // 'd1655
      11'd994  : in_data <= 14'h09a5; // 'd2469
      11'd995  : in_data <= 14'h153b; // 'd5435
      11'd996  : in_data <= 14'h03a4; // 'd932
      11'd997  : in_data <= 14'h1971; // 'd6513
      11'd998  : in_data <= 14'h1b3d; // 'd6973
      11'd999  : in_data <= 14'h0495; // 'd1173
      11'd1000 : in_data <= 14'h1b0e; // 'd6926
      11'd1001 : in_data <= 14'h0693; // 'd1683
      11'd1002 : in_data <= 14'h0517; // 'd1303
      11'd1003 : in_data <= 14'h1d6c; // 'd7532
      11'd1004 : in_data <= 14'h11e5; // 'd4581
      11'd1005 : in_data <= 14'h1bfc; // 'd7164
      11'd1006 : in_data <= 14'h069e; // 'd1694
      11'd1007 : in_data <= 14'h067b; // 'd1659
      11'd1008 : in_data <= 14'h096f; // 'd2415
      11'd1009 : in_data <= 14'h004b; // 'd75
      11'd1010 : in_data <= 14'h014a; // 'd330
      11'd1011 : in_data <= 14'h1926; // 'd6438
      11'd1012 : in_data <= 14'h141d; // 'd5149
      11'd1013 : in_data <= 14'h0148; // 'd328
      11'd1014 : in_data <= 14'h17b0; // 'd6064
      11'd1015 : in_data <= 14'h08db; // 'd2267
      11'd1016 : in_data <= 14'h16b9; // 'd5817
      11'd1017 : in_data <= 14'h1760; // 'd5984
      11'd1018 : in_data <= 14'h0825; // 'd2085
      11'd1019 : in_data <= 14'h0371; // 'd881
      11'd1020 : in_data <= 14'h14e1; // 'd5345
      11'd1021 : in_data <= 14'h0274; // 'd628
      11'd1022 : in_data <= 14'h0427; // 'd1063
      11'd1023 : in_data <= 14'h1852; // 'd6226
      11'd1024 : in_data <= 14'h18c0; // 'd6336
      11'd1025 : in_data <= 14'h06a4; // 'd1700
      11'd1026 : in_data <= 14'h11f7; // 'd4599
      11'd1027 : in_data <= 14'h0160; // 'd352
      11'd1028 : in_data <= 14'h0193; // 'd403
      11'd1029 : in_data <= 14'h088a; // 'd2186
      11'd1030 : in_data <= 14'h1bef; // 'd7151
      11'd1031 : in_data <= 14'h00a6; // 'd166
      11'd1032 : in_data <= 14'h1d95; // 'd7573
      11'd1033 : in_data <= 14'h0b75; // 'd2933
      11'd1034 : in_data <= 14'h0f1d; // 'd3869
      11'd1035 : in_data <= 14'h072e; // 'd1838
      11'd1036 : in_data <= 14'h050e; // 'd1294
      11'd1037 : in_data <= 14'h0f67; // 'd3943
      11'd1038 : in_data <= 14'h1731; // 'd5937
      11'd1039 : in_data <= 14'h0ec4; // 'd3780
      11'd1040 : in_data <= 14'h155c; // 'd5468
      11'd1041 : in_data <= 14'h0126; // 'd294
      11'd1042 : in_data <= 14'h0ce2; // 'd3298
      11'd1043 : in_data <= 14'h10d2; // 'd4306
      11'd1044 : in_data <= 14'h0a90; // 'd2704
      11'd1045 : in_data <= 14'h19a9; // 'd6569
      11'd1046 : in_data <= 14'h1061; // 'd4193
      11'd1047 : in_data <= 14'h0686; // 'd1670
      11'd1048 : in_data <= 14'h1758; // 'd5976
      11'd1049 : in_data <= 14'h04af; // 'd1199
      11'd1050 : in_data <= 14'h0369; // 'd873
      11'd1051 : in_data <= 14'h10e7; // 'd4327
      11'd1052 : in_data <= 14'h1499; // 'd5273
      11'd1053 : in_data <= 14'h11dc; // 'd4572
      11'd1054 : in_data <= 14'h13f2; // 'd5106
      11'd1055 : in_data <= 14'h1a2d; // 'd6701
      11'd1056 : in_data <= 14'h11ca; // 'd4554
      11'd1057 : in_data <= 14'h0a45; // 'd2629
      11'd1058 : in_data <= 14'h159c; // 'd5532
      11'd1059 : in_data <= 14'h14c5; // 'd5317
      11'd1060 : in_data <= 14'h060f; // 'd1551
      11'd1061 : in_data <= 14'h1387; // 'd4999
      11'd1062 : in_data <= 14'h1ae7; // 'd6887
      11'd1063 : in_data <= 14'h063c; // 'd1596
      11'd1064 : in_data <= 14'h1adf; // 'd6879
      11'd1065 : in_data <= 14'h10b1; // 'd4273
      11'd1066 : in_data <= 14'h19d5; // 'd6613
      11'd1067 : in_data <= 14'h05ef; // 'd1519
      11'd1068 : in_data <= 14'h044c; // 'd1100
      11'd1069 : in_data <= 14'h081f; // 'd2079
      11'd1070 : in_data <= 14'h0872; // 'd2162
      11'd1071 : in_data <= 14'h00dd; // 'd221
      11'd1072 : in_data <= 14'h1dc6; // 'd7622
      11'd1073 : in_data <= 14'h0d89; // 'd3465
      11'd1074 : in_data <= 14'h03fc; // 'd1020
      11'd1075 : in_data <= 14'h0c68; // 'd3176
      11'd1076 : in_data <= 14'h0742; // 'd1858
      11'd1077 : in_data <= 14'h03d3; // 'd979
      11'd1078 : in_data <= 14'h1440; // 'd5184
      11'd1079 : in_data <= 14'h0ebb; // 'd3771
      11'd1080 : in_data <= 14'h17b6; // 'd6070
      11'd1081 : in_data <= 14'h17be; // 'd6078
      11'd1082 : in_data <= 14'h09e5; // 'd2533
      11'd1083 : in_data <= 14'h1b3c; // 'd6972
      11'd1084 : in_data <= 14'h01cd; // 'd461
      11'd1085 : in_data <= 14'h0f8a; // 'd3978
      11'd1086 : in_data <= 14'h1471; // 'd5233
      11'd1087 : in_data <= 14'h032d; // 'd813
      11'd1088 : in_data <= 14'h1ec2; // 'd7874
      11'd1089 : in_data <= 14'h1ddd; // 'd7645
      11'd1090 : in_data <= 14'h0e88; // 'd3720
      11'd1091 : in_data <= 14'h0259; // 'd601
      11'd1092 : in_data <= 14'h09fd; // 'd2557
      11'd1093 : in_data <= 14'h16bc; // 'd5820
      11'd1094 : in_data <= 14'h102f; // 'd4143
      11'd1095 : in_data <= 14'h1bb9; // 'd7097
      11'd1096 : in_data <= 14'h13a0; // 'd5024
      11'd1097 : in_data <= 14'h04bd; // 'd1213
      11'd1098 : in_data <= 14'h1d9c; // 'd7580
      11'd1099 : in_data <= 14'h1ec2; // 'd7874
      11'd1100 : in_data <= 14'h04e9; // 'd1257
      11'd1101 : in_data <= 14'h1a6d; // 'd6765
      11'd1102 : in_data <= 14'h165e; // 'd5726
      11'd1103 : in_data <= 14'h10a9; // 'd4265
      11'd1104 : in_data <= 14'h19c0; // 'd6592
      11'd1105 : in_data <= 14'h03b7; // 'd951
      11'd1106 : in_data <= 14'h1483; // 'd5251
      11'd1107 : in_data <= 14'h09a3; // 'd2467
      11'd1108 : in_data <= 14'h0e73; // 'd3699
      11'd1109 : in_data <= 14'h1a9f; // 'd6815
      11'd1110 : in_data <= 14'h0407; // 'd1031
      11'd1111 : in_data <= 14'h028c; // 'd652
      11'd1112 : in_data <= 14'h1e26; // 'd7718
      11'd1113 : in_data <= 14'h0996; // 'd2454
      11'd1114 : in_data <= 14'h0d9c; // 'd3484
      11'd1115 : in_data <= 14'h0397; // 'd919
      11'd1116 : in_data <= 14'h01f3; // 'd499
      11'd1117 : in_data <= 14'h1467; // 'd5223
      11'd1118 : in_data <= 14'h145c; // 'd5212
      11'd1119 : in_data <= 14'h1a0a; // 'd6666
      11'd1120 : in_data <= 14'h0472; // 'd1138
      11'd1121 : in_data <= 14'h065c; // 'd1628
      11'd1122 : in_data <= 14'h0b0d; // 'd2829
      11'd1123 : in_data <= 14'h03e6; // 'd998
      11'd1124 : in_data <= 14'h0e64; // 'd3684
      11'd1125 : in_data <= 14'h121a; // 'd4634
      11'd1126 : in_data <= 14'h1d6e; // 'd7534
      11'd1127 : in_data <= 14'h0679; // 'd1657
      11'd1128 : in_data <= 14'h1c34; // 'd7220
      11'd1129 : in_data <= 14'h1d8f; // 'd7567
      11'd1130 : in_data <= 14'h01cf; // 'd463
      11'd1131 : in_data <= 14'h17dc; // 'd6108
      11'd1132 : in_data <= 14'h1b97; // 'd7063
      11'd1133 : in_data <= 14'h04f8; // 'd1272
      11'd1134 : in_data <= 14'h1684; // 'd5764
      11'd1135 : in_data <= 14'h1b2d; // 'd6957
      11'd1136 : in_data <= 14'h05ed; // 'd1517
      11'd1137 : in_data <= 14'h1ba9; // 'd7081
      11'd1138 : in_data <= 14'h0332; // 'd818
      11'd1139 : in_data <= 14'h04e8; // 'd1256
      11'd1140 : in_data <= 14'h1c3a; // 'd7226
      11'd1141 : in_data <= 14'h1258; // 'd4696
      11'd1142 : in_data <= 14'h1c16; // 'd7190
      11'd1143 : in_data <= 14'h0f1d; // 'd3869
      11'd1144 : in_data <= 14'h06f9; // 'd1785
      11'd1145 : in_data <= 14'h1a14; // 'd6676
      11'd1146 : in_data <= 14'h00f9; // 'd249
      11'd1147 : in_data <= 14'h173c; // 'd5948
      11'd1148 : in_data <= 14'h1d9b; // 'd7579
      11'd1149 : in_data <= 14'h0941; // 'd2369
      11'd1150 : in_data <= 14'h013b; // 'd315
      11'd1151 : in_data <= 14'h12a2; // 'd4770
      11'd1152 : in_data <= 14'h1478; // 'd5240
      11'd1153 : in_data <= 14'h16e2; // 'd5858
      11'd1154 : in_data <= 14'h0f02; // 'd3842
      11'd1155 : in_data <= 14'h0232; // 'd562
      11'd1156 : in_data <= 14'h0239; // 'd569
      11'd1157 : in_data <= 14'h0bc0; // 'd3008
      11'd1158 : in_data <= 14'h0705; // 'd1797
      11'd1159 : in_data <= 14'h0bd2; // 'd3026
      11'd1160 : in_data <= 14'h1cda; // 'd7386
      11'd1161 : in_data <= 14'h0b1b; // 'd2843
      11'd1162 : in_data <= 14'h162f; // 'd5679
      11'd1163 : in_data <= 14'h1287; // 'd4743
      11'd1164 : in_data <= 14'h1c57; // 'd7255
      11'd1165 : in_data <= 14'h1bd5; // 'd7125
      11'd1166 : in_data <= 14'h1d33; // 'd7475
      11'd1167 : in_data <= 14'h1d9a; // 'd7578
      11'd1168 : in_data <= 14'h1ad0; // 'd6864
      11'd1169 : in_data <= 14'h1bdf; // 'd7135
      11'd1170 : in_data <= 14'h148d; // 'd5261
      11'd1171 : in_data <= 14'h06f1; // 'd1777
      11'd1172 : in_data <= 14'h0cd4; // 'd3284
      11'd1173 : in_data <= 14'h15bd; // 'd5565
      11'd1174 : in_data <= 14'h14e4; // 'd5348
      11'd1175 : in_data <= 14'h071d; // 'd1821
      11'd1176 : in_data <= 14'h1c87; // 'd7303
      11'd1177 : in_data <= 14'h1264; // 'd4708
      11'd1178 : in_data <= 14'h149d; // 'd5277
      11'd1179 : in_data <= 14'h0c12; // 'd3090
      11'd1180 : in_data <= 14'h0841; // 'd2113
      11'd1181 : in_data <= 14'h1166; // 'd4454
      11'd1182 : in_data <= 14'h087f; // 'd2175
      11'd1183 : in_data <= 14'h0c7f; // 'd3199
      11'd1184 : in_data <= 14'h000e; // 'd14
      11'd1185 : in_data <= 14'h1d30; // 'd7472
      11'd1186 : in_data <= 14'h1c8a; // 'd7306
      11'd1187 : in_data <= 14'h1ba9; // 'd7081
      11'd1188 : in_data <= 14'h151c; // 'd5404
      11'd1189 : in_data <= 14'h1e10; // 'd7696
      11'd1190 : in_data <= 14'h0015; // 'd21
      11'd1191 : in_data <= 14'h0773; // 'd1907
      11'd1192 : in_data <= 14'h1a03; // 'd6659
      11'd1193 : in_data <= 14'h0714; // 'd1812
      11'd1194 : in_data <= 14'h19e8; // 'd6632
      11'd1195 : in_data <= 14'h0148; // 'd328
      11'd1196 : in_data <= 14'h11da; // 'd4570
      11'd1197 : in_data <= 14'h1de9; // 'd7657
      11'd1198 : in_data <= 14'h1b31; // 'd6961
      11'd1199 : in_data <= 14'h1a96; // 'd6806
      11'd1200 : in_data <= 14'h116b; // 'd4459
      11'd1201 : in_data <= 14'h19b1; // 'd6577
      11'd1202 : in_data <= 14'h0287; // 'd647
      11'd1203 : in_data <= 14'h01ac; // 'd428
      11'd1204 : in_data <= 14'h1908; // 'd6408
      11'd1205 : in_data <= 14'h047c; // 'd1148
      11'd1206 : in_data <= 14'h0a8e; // 'd2702
      11'd1207 : in_data <= 14'h0aad; // 'd2733
      11'd1208 : in_data <= 14'h14a9; // 'd5289
      11'd1209 : in_data <= 14'h1cc4; // 'd7364
      11'd1210 : in_data <= 14'h115c; // 'd4444
      11'd1211 : in_data <= 14'h1a89; // 'd6793
      11'd1212 : in_data <= 14'h08a6; // 'd2214
      11'd1213 : in_data <= 14'h0b26; // 'd2854
      11'd1214 : in_data <= 14'h1617; // 'd5655
      11'd1215 : in_data <= 14'h0d0b; // 'd3339
      11'd1216 : in_data <= 14'h1120; // 'd4384
      11'd1217 : in_data <= 14'h049c; // 'd1180
      11'd1218 : in_data <= 14'h0622; // 'd1570
      11'd1219 : in_data <= 14'h10d5; // 'd4309
      11'd1220 : in_data <= 14'h1477; // 'd5239
      11'd1221 : in_data <= 14'h1cc4; // 'd7364
      11'd1222 : in_data <= 14'h1546; // 'd5446
      11'd1223 : in_data <= 14'h07c1; // 'd1985
      11'd1224 : in_data <= 14'h0541; // 'd1345
      11'd1225 : in_data <= 14'h18ee; // 'd6382
      11'd1226 : in_data <= 14'h049a; // 'd1178
      11'd1227 : in_data <= 14'h0648; // 'd1608
      11'd1228 : in_data <= 14'h16e8; // 'd5864
      11'd1229 : in_data <= 14'h07c5; // 'd1989
      11'd1230 : in_data <= 14'h067d; // 'd1661
      11'd1231 : in_data <= 14'h1c05; // 'd7173
      11'd1232 : in_data <= 14'h0bf1; // 'd3057
      11'd1233 : in_data <= 14'h04fa; // 'd1274
      11'd1234 : in_data <= 14'h171c; // 'd5916
      11'd1235 : in_data <= 14'h0d62; // 'd3426
      11'd1236 : in_data <= 14'h0b7b; // 'd2939
      11'd1237 : in_data <= 14'h065a; // 'd1626
      11'd1238 : in_data <= 14'h066e; // 'd1646
      11'd1239 : in_data <= 14'h1e8f; // 'd7823
      11'd1240 : in_data <= 14'h1a4b; // 'd6731
      11'd1241 : in_data <= 14'h083c; // 'd2108
      11'd1242 : in_data <= 14'h16ee; // 'd5870
      11'd1243 : in_data <= 14'h0eef; // 'd3823
      11'd1244 : in_data <= 14'h14b9; // 'd5305
      11'd1245 : in_data <= 14'h076a; // 'd1898
      11'd1246 : in_data <= 14'h0e18; // 'd3608
      11'd1247 : in_data <= 14'h0e5b; // 'd3675
      11'd1248 : in_data <= 14'h01ab; // 'd427
      11'd1249 : in_data <= 14'h19c8; // 'd6600
      11'd1250 : in_data <= 14'h1298; // 'd4760
      11'd1251 : in_data <= 14'h1975; // 'd6517
      11'd1252 : in_data <= 14'h0b26; // 'd2854
      11'd1253 : in_data <= 14'h048a; // 'd1162
      11'd1254 : in_data <= 14'h1883; // 'd6275
      11'd1255 : in_data <= 14'h1a90; // 'd6800
      11'd1256 : in_data <= 14'h0d1e; // 'd3358
      11'd1257 : in_data <= 14'h1db5; // 'd7605
      11'd1258 : in_data <= 14'h0978; // 'd2424
      11'd1259 : in_data <= 14'h1529; // 'd5417
      11'd1260 : in_data <= 14'h0df0; // 'd3568
      11'd1261 : in_data <= 14'h015b; // 'd347
      11'd1262 : in_data <= 14'h01d2; // 'd466
      11'd1263 : in_data <= 14'h0bae; // 'd2990
      11'd1264 : in_data <= 14'h1ebc; // 'd7868
      11'd1265 : in_data <= 14'h12a2; // 'd4770
      11'd1266 : in_data <= 14'h0f1e; // 'd3870
      11'd1267 : in_data <= 14'h0688; // 'd1672
      11'd1268 : in_data <= 14'h071a; // 'd1818
      11'd1269 : in_data <= 14'h0722; // 'd1826
      11'd1270 : in_data <= 14'h0828; // 'd2088
      11'd1271 : in_data <= 14'h12b1; // 'd4785
      11'd1272 : in_data <= 14'h1120; // 'd4384
      11'd1273 : in_data <= 14'h00a7; // 'd167
      11'd1274 : in_data <= 14'h1270; // 'd4720
      11'd1275 : in_data <= 14'h1d01; // 'd7425
      11'd1276 : in_data <= 14'h16ec; // 'd5868
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      12'd0    : out_data_ref <= 8'h52;
      12'd1    : out_data_ref <= 8'hb4;
      12'd2    : out_data_ref <= 8'h1f;
      12'd3    : out_data_ref <= 8'h04;
      12'd4    : out_data_ref <= 8'hf8;
      12'd5    : out_data_ref <= 8'h3b;
      12'd6    : out_data_ref <= 8'h7e;
      12'd7    : out_data_ref <= 8'hba;
      12'd8    : out_data_ref <= 8'h97;
      12'd9    : out_data_ref <= 8'hb1;
      12'd10   : out_data_ref <= 8'h9f;
      12'd11   : out_data_ref <= 8'ha0;
      12'd12   : out_data_ref <= 8'h5e;
      12'd13   : out_data_ref <= 8'h55;
      12'd14   : out_data_ref <= 8'h22;
      12'd15   : out_data_ref <= 8'he9;
      12'd16   : out_data_ref <= 8'he8;
      12'd17   : out_data_ref <= 8'hed;
      12'd18   : out_data_ref <= 8'hde;
      12'd19   : out_data_ref <= 8'h6a;
      12'd20   : out_data_ref <= 8'h15;
      12'd21   : out_data_ref <= 8'h0d;
      12'd22   : out_data_ref <= 8'hfd;
      12'd23   : out_data_ref <= 8'he7;
      12'd24   : out_data_ref <= 8'hdc;
      12'd25   : out_data_ref <= 8'hb9;
      12'd26   : out_data_ref <= 8'he9;
      12'd27   : out_data_ref <= 8'h01;
      12'd28   : out_data_ref <= 8'hf4;
      12'd29   : out_data_ref <= 8'h8b;
      12'd30   : out_data_ref <= 8'h76;
      12'd31   : out_data_ref <= 8'h30;
      12'd32   : out_data_ref <= 8'h83;
      12'd33   : out_data_ref <= 8'h60;
      12'd34   : out_data_ref <= 8'h7a;
      12'd35   : out_data_ref <= 8'hfc;
      12'd36   : out_data_ref <= 8'h0b;
      12'd37   : out_data_ref <= 8'h35;
      12'd38   : out_data_ref <= 8'ha7;
      12'd39   : out_data_ref <= 8'h80;
      12'd40   : out_data_ref <= 8'he0;
      12'd41   : out_data_ref <= 8'h96;
      12'd42   : out_data_ref <= 8'hea;
      12'd43   : out_data_ref <= 8'hbe;
      12'd44   : out_data_ref <= 8'ha9;
      12'd45   : out_data_ref <= 8'h88;
      12'd46   : out_data_ref <= 8'h1e;
      12'd47   : out_data_ref <= 8'hd0;
      12'd48   : out_data_ref <= 8'hae;
      12'd49   : out_data_ref <= 8'hfd;
      12'd50   : out_data_ref <= 8'h75;
      12'd51   : out_data_ref <= 8'h35;
      12'd52   : out_data_ref <= 8'h83;
      12'd53   : out_data_ref <= 8'h84;
      12'd54   : out_data_ref <= 8'h39;
      12'd55   : out_data_ref <= 8'h28;
      12'd56   : out_data_ref <= 8'h0d;
      12'd57   : out_data_ref <= 8'hf3;
      12'd58   : out_data_ref <= 8'h5d;
      12'd59   : out_data_ref <= 8'h77;
      12'd60   : out_data_ref <= 8'h8b;
      12'd61   : out_data_ref <= 8'h98;
      12'd62   : out_data_ref <= 8'h89;
      12'd63   : out_data_ref <= 8'hce;
      12'd64   : out_data_ref <= 8'h25;
      12'd65   : out_data_ref <= 8'h08;
      12'd66   : out_data_ref <= 8'h4b;
      12'd67   : out_data_ref <= 8'hd1;
      12'd68   : out_data_ref <= 8'h7a;
      12'd69   : out_data_ref <= 8'hb5;
      12'd70   : out_data_ref <= 8'h1e;
      12'd71   : out_data_ref <= 8'hd8;
      12'd72   : out_data_ref <= 8'hde;
      12'd73   : out_data_ref <= 8'h60;
      12'd74   : out_data_ref <= 8'h33;
      12'd75   : out_data_ref <= 8'h71;
      12'd76   : out_data_ref <= 8'h76;
      12'd77   : out_data_ref <= 8'h5f;
      12'd78   : out_data_ref <= 8'h5c;
      12'd79   : out_data_ref <= 8'hc9;
      12'd80   : out_data_ref <= 8'hba;
      12'd81   : out_data_ref <= 8'h4b;
      12'd82   : out_data_ref <= 8'h3e;
      12'd83   : out_data_ref <= 8'h03;
      12'd84   : out_data_ref <= 8'hc9;
      12'd85   : out_data_ref <= 8'h0f;
      12'd86   : out_data_ref <= 8'h83;
      12'd87   : out_data_ref <= 8'h95;
      12'd88   : out_data_ref <= 8'h0d;
      12'd89   : out_data_ref <= 8'h7b;
      12'd90   : out_data_ref <= 8'h82;
      12'd91   : out_data_ref <= 8'h8e;
      12'd92   : out_data_ref <= 8'h2e;
      12'd93   : out_data_ref <= 8'h3e;
      12'd94   : out_data_ref <= 8'hc7;
      12'd95   : out_data_ref <= 8'h0a;
      12'd96   : out_data_ref <= 8'h7f;
      12'd97   : out_data_ref <= 8'h2b;
      12'd98   : out_data_ref <= 8'h87;
      12'd99   : out_data_ref <= 8'h5e;
      12'd100  : out_data_ref <= 8'hd3;
      12'd101  : out_data_ref <= 8'h8a;
      12'd102  : out_data_ref <= 8'h70;
      12'd103  : out_data_ref <= 8'hac;
      12'd104  : out_data_ref <= 8'h4a;
      12'd105  : out_data_ref <= 8'h81;
      12'd106  : out_data_ref <= 8'h26;
      12'd107  : out_data_ref <= 8'h32;
      12'd108  : out_data_ref <= 8'h7a;
      12'd109  : out_data_ref <= 8'hc2;
      12'd110  : out_data_ref <= 8'hc0;
      12'd111  : out_data_ref <= 8'hd2;
      12'd112  : out_data_ref <= 8'hb4;
      12'd113  : out_data_ref <= 8'h61;
      12'd114  : out_data_ref <= 8'h99;
      12'd115  : out_data_ref <= 8'h9a;
      12'd116  : out_data_ref <= 8'h81;
      12'd117  : out_data_ref <= 8'h30;
      12'd118  : out_data_ref <= 8'hd1;
      12'd119  : out_data_ref <= 8'hef;
      12'd120  : out_data_ref <= 8'h2f;
      12'd121  : out_data_ref <= 8'hb7;
      12'd122  : out_data_ref <= 8'h50;
      12'd123  : out_data_ref <= 8'h2d;
      12'd124  : out_data_ref <= 8'h29;
      12'd125  : out_data_ref <= 8'hbc;
      12'd126  : out_data_ref <= 8'h33;
      12'd127  : out_data_ref <= 8'h75;
      12'd128  : out_data_ref <= 8'h22;
      12'd129  : out_data_ref <= 8'h39;
      12'd130  : out_data_ref <= 8'hca;
      12'd131  : out_data_ref <= 8'h3e;
      12'd132  : out_data_ref <= 8'h64;
      12'd133  : out_data_ref <= 8'h17;
      12'd134  : out_data_ref <= 8'h53;
      12'd135  : out_data_ref <= 8'h7c;
      12'd136  : out_data_ref <= 8'h6c;
      12'd137  : out_data_ref <= 8'h2b;
      12'd138  : out_data_ref <= 8'h03;
      12'd139  : out_data_ref <= 8'h91;
      12'd140  : out_data_ref <= 8'h51;
      12'd141  : out_data_ref <= 8'h45;
      12'd142  : out_data_ref <= 8'hdd;
      12'd143  : out_data_ref <= 8'h7d;
      12'd144  : out_data_ref <= 8'ha8;
      12'd145  : out_data_ref <= 8'h00;
      12'd146  : out_data_ref <= 8'h2b;
      12'd147  : out_data_ref <= 8'h35;
      12'd148  : out_data_ref <= 8'haa;
      12'd149  : out_data_ref <= 8'h9a;
      12'd150  : out_data_ref <= 8'h90;
      12'd151  : out_data_ref <= 8'haa;
      12'd152  : out_data_ref <= 8'h08;
      12'd153  : out_data_ref <= 8'h27;
      12'd154  : out_data_ref <= 8'h53;
      12'd155  : out_data_ref <= 8'h3c;
      12'd156  : out_data_ref <= 8'h51;
      12'd157  : out_data_ref <= 8'h7a;
      12'd158  : out_data_ref <= 8'hc3;
      12'd159  : out_data_ref <= 8'h73;
      12'd160  : out_data_ref <= 8'hc0;
      12'd161  : out_data_ref <= 8'ha8;
      12'd162  : out_data_ref <= 8'hd6;
      12'd163  : out_data_ref <= 8'hfa;
      12'd164  : out_data_ref <= 8'h51;
      12'd165  : out_data_ref <= 8'h9d;
      12'd166  : out_data_ref <= 8'h9a;
      12'd167  : out_data_ref <= 8'h77;
      12'd168  : out_data_ref <= 8'hd5;
      12'd169  : out_data_ref <= 8'h6b;
      12'd170  : out_data_ref <= 8'h2a;
      12'd171  : out_data_ref <= 8'hca;
      12'd172  : out_data_ref <= 8'ha0;
      12'd173  : out_data_ref <= 8'h9b;
      12'd174  : out_data_ref <= 8'ha7;
      12'd175  : out_data_ref <= 8'h01;
      12'd176  : out_data_ref <= 8'hbc;
      12'd177  : out_data_ref <= 8'h18;
      12'd178  : out_data_ref <= 8'h1c;
      12'd179  : out_data_ref <= 8'hb1;
      12'd180  : out_data_ref <= 8'h67;
      12'd181  : out_data_ref <= 8'hf8;
      12'd182  : out_data_ref <= 8'hf1;
      12'd183  : out_data_ref <= 8'hc0;
      12'd184  : out_data_ref <= 8'hfe;
      12'd185  : out_data_ref <= 8'ha5;
      12'd186  : out_data_ref <= 8'h2d;
      12'd187  : out_data_ref <= 8'h45;
      12'd188  : out_data_ref <= 8'had;
      12'd189  : out_data_ref <= 8'hec;
      12'd190  : out_data_ref <= 8'h44;
      12'd191  : out_data_ref <= 8'hbe;
      12'd192  : out_data_ref <= 8'hc9;
      12'd193  : out_data_ref <= 8'h38;
      12'd194  : out_data_ref <= 8'h85;
      12'd195  : out_data_ref <= 8'h85;
      12'd196  : out_data_ref <= 8'hae;
      12'd197  : out_data_ref <= 8'hcb;
      12'd198  : out_data_ref <= 8'ha6;
      12'd199  : out_data_ref <= 8'h1e;
      12'd200  : out_data_ref <= 8'hd3;
      12'd201  : out_data_ref <= 8'h13;
      12'd202  : out_data_ref <= 8'h0d;
      12'd203  : out_data_ref <= 8'h09;
      12'd204  : out_data_ref <= 8'h99;
      12'd205  : out_data_ref <= 8'hc5;
      12'd206  : out_data_ref <= 8'h43;
      12'd207  : out_data_ref <= 8'h0f;
      12'd208  : out_data_ref <= 8'hc0;
      12'd209  : out_data_ref <= 8'hee;
      12'd210  : out_data_ref <= 8'h79;
      12'd211  : out_data_ref <= 8'h0a;
      12'd212  : out_data_ref <= 8'h4c;
      12'd213  : out_data_ref <= 8'hcd;
      12'd214  : out_data_ref <= 8'h73;
      12'd215  : out_data_ref <= 8'h5e;
      12'd216  : out_data_ref <= 8'hf3;
      12'd217  : out_data_ref <= 8'h84;
      12'd218  : out_data_ref <= 8'hd2;
      12'd219  : out_data_ref <= 8'hc5;
      12'd220  : out_data_ref <= 8'hcd;
      12'd221  : out_data_ref <= 8'h90;
      12'd222  : out_data_ref <= 8'h48;
      12'd223  : out_data_ref <= 8'hb5;
      12'd224  : out_data_ref <= 8'h4f;
      12'd225  : out_data_ref <= 8'he7;
      12'd226  : out_data_ref <= 8'h75;
      12'd227  : out_data_ref <= 8'h78;
      12'd228  : out_data_ref <= 8'hba;
      12'd229  : out_data_ref <= 8'h3e;
      12'd230  : out_data_ref <= 8'hfb;
      12'd231  : out_data_ref <= 8'hcb;
      12'd232  : out_data_ref <= 8'h51;
      12'd233  : out_data_ref <= 8'hef;
      12'd234  : out_data_ref <= 8'h5d;
      12'd235  : out_data_ref <= 8'ha2;
      12'd236  : out_data_ref <= 8'h2b;
      12'd237  : out_data_ref <= 8'hea;
      12'd238  : out_data_ref <= 8'hca;
      12'd239  : out_data_ref <= 8'h98;
      12'd240  : out_data_ref <= 8'h97;
      12'd241  : out_data_ref <= 8'h79;
      12'd242  : out_data_ref <= 8'hfe;
      12'd243  : out_data_ref <= 8'h47;
      12'd244  : out_data_ref <= 8'he8;
      12'd245  : out_data_ref <= 8'h97;
      12'd246  : out_data_ref <= 8'h92;
      12'd247  : out_data_ref <= 8'h41;
      12'd248  : out_data_ref <= 8'h60;
      12'd249  : out_data_ref <= 8'hca;
      12'd250  : out_data_ref <= 8'h37;
      12'd251  : out_data_ref <= 8'h34;
      12'd252  : out_data_ref <= 8'hcb;
      12'd253  : out_data_ref <= 8'h3f;
      12'd254  : out_data_ref <= 8'hfa;
      12'd255  : out_data_ref <= 8'h07;
      12'd256  : out_data_ref <= 8'h5f;
      12'd257  : out_data_ref <= 8'h29;
      12'd258  : out_data_ref <= 8'h49;
      12'd259  : out_data_ref <= 8'hee;
      12'd260  : out_data_ref <= 8'h23;
      12'd261  : out_data_ref <= 8'h69;
      12'd262  : out_data_ref <= 8'ha0;
      12'd263  : out_data_ref <= 8'hb0;
      12'd264  : out_data_ref <= 8'hc7;
      12'd265  : out_data_ref <= 8'h9d;
      12'd266  : out_data_ref <= 8'he5;
      12'd267  : out_data_ref <= 8'h0e;
      12'd268  : out_data_ref <= 8'h0d;
      12'd269  : out_data_ref <= 8'h2b;
      12'd270  : out_data_ref <= 8'hca;
      12'd271  : out_data_ref <= 8'h0a;
      12'd272  : out_data_ref <= 8'hd6;
      12'd273  : out_data_ref <= 8'h95;
      12'd274  : out_data_ref <= 8'h3a;
      12'd275  : out_data_ref <= 8'h71;
      12'd276  : out_data_ref <= 8'h97;
      12'd277  : out_data_ref <= 8'hcd;
      12'd278  : out_data_ref <= 8'h23;
      12'd279  : out_data_ref <= 8'h19;
      12'd280  : out_data_ref <= 8'hfd;
      12'd281  : out_data_ref <= 8'h68;
      12'd282  : out_data_ref <= 8'h19;
      12'd283  : out_data_ref <= 8'hec;
      12'd284  : out_data_ref <= 8'h25;
      12'd285  : out_data_ref <= 8'ha9;
      12'd286  : out_data_ref <= 8'h1c;
      12'd287  : out_data_ref <= 8'h37;
      12'd288  : out_data_ref <= 8'h6b;
      12'd289  : out_data_ref <= 8'h83;
      12'd290  : out_data_ref <= 8'h14;
      12'd291  : out_data_ref <= 8'hd9;
      12'd292  : out_data_ref <= 8'h25;
      12'd293  : out_data_ref <= 8'h23;
      12'd294  : out_data_ref <= 8'hc7;
      12'd295  : out_data_ref <= 8'haa;
      12'd296  : out_data_ref <= 8'ha6;
      12'd297  : out_data_ref <= 8'h01;
      12'd298  : out_data_ref <= 8'h4f;
      12'd299  : out_data_ref <= 8'hdc;
      12'd300  : out_data_ref <= 8'h0d;
      12'd301  : out_data_ref <= 8'h45;
      12'd302  : out_data_ref <= 8'h3b;
      12'd303  : out_data_ref <= 8'h6a;
      12'd304  : out_data_ref <= 8'h81;
      12'd305  : out_data_ref <= 8'h4e;
      12'd306  : out_data_ref <= 8'ha7;
      12'd307  : out_data_ref <= 8'h15;
      12'd308  : out_data_ref <= 8'h3f;
      12'd309  : out_data_ref <= 8'h82;
      12'd310  : out_data_ref <= 8'h7d;
      12'd311  : out_data_ref <= 8'he0;
      12'd312  : out_data_ref <= 8'h3f;
      12'd313  : out_data_ref <= 8'h47;
      12'd314  : out_data_ref <= 8'h0a;
      12'd315  : out_data_ref <= 8'h10;
      12'd316  : out_data_ref <= 8'hde;
      12'd317  : out_data_ref <= 8'ha5;
      12'd318  : out_data_ref <= 8'h22;
      12'd319  : out_data_ref <= 8'h6b;
      12'd320  : out_data_ref <= 8'hfb;
      12'd321  : out_data_ref <= 8'hb2;
      12'd322  : out_data_ref <= 8'hca;
      12'd323  : out_data_ref <= 8'hcd;
      12'd324  : out_data_ref <= 8'h41;
      12'd325  : out_data_ref <= 8'heb;
      12'd326  : out_data_ref <= 8'hec;
      12'd327  : out_data_ref <= 8'haa;
      12'd328  : out_data_ref <= 8'h8c;
      12'd329  : out_data_ref <= 8'h84;
      12'd330  : out_data_ref <= 8'hbc;
      12'd331  : out_data_ref <= 8'h19;
      12'd332  : out_data_ref <= 8'h38;
      12'd333  : out_data_ref <= 8'hd8;
      12'd334  : out_data_ref <= 8'h03;
      12'd335  : out_data_ref <= 8'h9b;
      12'd336  : out_data_ref <= 8'h06;
      12'd337  : out_data_ref <= 8'h68;
      12'd338  : out_data_ref <= 8'h74;
      12'd339  : out_data_ref <= 8'h7a;
      12'd340  : out_data_ref <= 8'h99;
      12'd341  : out_data_ref <= 8'h9f;
      12'd342  : out_data_ref <= 8'h90;
      12'd343  : out_data_ref <= 8'he2;
      12'd344  : out_data_ref <= 8'h9c;
      12'd345  : out_data_ref <= 8'h22;
      12'd346  : out_data_ref <= 8'hca;
      12'd347  : out_data_ref <= 8'had;
      12'd348  : out_data_ref <= 8'h88;
      12'd349  : out_data_ref <= 8'h91;
      12'd350  : out_data_ref <= 8'h8f;
      12'd351  : out_data_ref <= 8'h22;
      12'd352  : out_data_ref <= 8'h16;
      12'd353  : out_data_ref <= 8'h6a;
      12'd354  : out_data_ref <= 8'h9f;
      12'd355  : out_data_ref <= 8'h97;
      12'd356  : out_data_ref <= 8'he8;
      12'd357  : out_data_ref <= 8'hc8;
      12'd358  : out_data_ref <= 8'h2c;
      12'd359  : out_data_ref <= 8'hc9;
      12'd360  : out_data_ref <= 8'hbe;
      12'd361  : out_data_ref <= 8'he1;
      12'd362  : out_data_ref <= 8'hef;
      12'd363  : out_data_ref <= 8'hf6;
      12'd364  : out_data_ref <= 8'hb3;
      12'd365  : out_data_ref <= 8'hbb;
      12'd366  : out_data_ref <= 8'ha8;
      12'd367  : out_data_ref <= 8'hb7;
      12'd368  : out_data_ref <= 8'he3;
      12'd369  : out_data_ref <= 8'hd0;
      12'd370  : out_data_ref <= 8'h5c;
      12'd371  : out_data_ref <= 8'hbc;
      12'd372  : out_data_ref <= 8'h8d;
      12'd373  : out_data_ref <= 8'h26;
      12'd374  : out_data_ref <= 8'ha3;
      12'd375  : out_data_ref <= 8'h64;
      12'd376  : out_data_ref <= 8'h45;
      12'd377  : out_data_ref <= 8'h0d;
      12'd378  : out_data_ref <= 8'h43;
      12'd379  : out_data_ref <= 8'hf8;
      12'd380  : out_data_ref <= 8'h56;
      12'd381  : out_data_ref <= 8'h1a;
      12'd382  : out_data_ref <= 8'h5a;
      12'd383  : out_data_ref <= 8'h59;
      12'd384  : out_data_ref <= 8'h8c;
      12'd385  : out_data_ref <= 8'h69;
      12'd386  : out_data_ref <= 8'hac;
      12'd387  : out_data_ref <= 8'h28;
      12'd388  : out_data_ref <= 8'hd5;
      12'd389  : out_data_ref <= 8'h34;
      12'd390  : out_data_ref <= 8'hf7;
      12'd391  : out_data_ref <= 8'hdd;
      12'd392  : out_data_ref <= 8'h4c;
      12'd393  : out_data_ref <= 8'h92;
      12'd394  : out_data_ref <= 8'hc2;
      12'd395  : out_data_ref <= 8'hdd;
      12'd396  : out_data_ref <= 8'he5;
      12'd397  : out_data_ref <= 8'hbe;
      12'd398  : out_data_ref <= 8'hb1;
      12'd399  : out_data_ref <= 8'hc6;
      12'd400  : out_data_ref <= 8'h4c;
      12'd401  : out_data_ref <= 8'h55;
      12'd402  : out_data_ref <= 8'ha7;
      12'd403  : out_data_ref <= 8'h32;
      12'd404  : out_data_ref <= 8'hb7;
      12'd405  : out_data_ref <= 8'h4e;
      12'd406  : out_data_ref <= 8'h9b;
      12'd407  : out_data_ref <= 8'h89;
      12'd408  : out_data_ref <= 8'h22;
      12'd409  : out_data_ref <= 8'h1d;
      12'd410  : out_data_ref <= 8'hb3;
      12'd411  : out_data_ref <= 8'h03;
      12'd412  : out_data_ref <= 8'h20;
      12'd413  : out_data_ref <= 8'hc7;
      12'd414  : out_data_ref <= 8'h71;
      12'd415  : out_data_ref <= 8'h99;
      12'd416  : out_data_ref <= 8'hf5;
      12'd417  : out_data_ref <= 8'h2b;
      12'd418  : out_data_ref <= 8'h08;
      12'd419  : out_data_ref <= 8'ha2;
      12'd420  : out_data_ref <= 8'h7b;
      12'd421  : out_data_ref <= 8'h7c;
      12'd422  : out_data_ref <= 8'hf3;
      12'd423  : out_data_ref <= 8'h43;
      12'd424  : out_data_ref <= 8'h7a;
      12'd425  : out_data_ref <= 8'h10;
      12'd426  : out_data_ref <= 8'hf5;
      12'd427  : out_data_ref <= 8'hb7;
      12'd428  : out_data_ref <= 8'h7c;
      12'd429  : out_data_ref <= 8'hbd;
      12'd430  : out_data_ref <= 8'h09;
      12'd431  : out_data_ref <= 8'h30;
      12'd432  : out_data_ref <= 8'hb0;
      12'd433  : out_data_ref <= 8'hbf;
      12'd434  : out_data_ref <= 8'hd8;
      12'd435  : out_data_ref <= 8'h46;
      12'd436  : out_data_ref <= 8'h28;
      12'd437  : out_data_ref <= 8'hcd;
      12'd438  : out_data_ref <= 8'hd1;
      12'd439  : out_data_ref <= 8'h29;
      12'd440  : out_data_ref <= 8'hd9;
      12'd441  : out_data_ref <= 8'hcf;
      12'd442  : out_data_ref <= 8'h9b;
      12'd443  : out_data_ref <= 8'heb;
      12'd444  : out_data_ref <= 8'hb9;
      12'd445  : out_data_ref <= 8'hca;
      12'd446  : out_data_ref <= 8'he0;
      12'd447  : out_data_ref <= 8'hc4;
      12'd448  : out_data_ref <= 8'hb4;
      12'd449  : out_data_ref <= 8'h14;
      12'd450  : out_data_ref <= 8'h91;
      12'd451  : out_data_ref <= 8'hd0;
      12'd452  : out_data_ref <= 8'h40;
      12'd453  : out_data_ref <= 8'h2f;
      12'd454  : out_data_ref <= 8'hf1;
      12'd455  : out_data_ref <= 8'h56;
      12'd456  : out_data_ref <= 8'h7a;
      12'd457  : out_data_ref <= 8'hf3;
      12'd458  : out_data_ref <= 8'h5b;
      12'd459  : out_data_ref <= 8'ha5;
      12'd460  : out_data_ref <= 8'h98;
      12'd461  : out_data_ref <= 8'hf2;
      12'd462  : out_data_ref <= 8'h9f;
      12'd463  : out_data_ref <= 8'hab;
      12'd464  : out_data_ref <= 8'hce;
      12'd465  : out_data_ref <= 8'h96;
      12'd466  : out_data_ref <= 8'had;
      12'd467  : out_data_ref <= 8'h8b;
      12'd468  : out_data_ref <= 8'h68;
      12'd469  : out_data_ref <= 8'hea;
      12'd470  : out_data_ref <= 8'h6f;
      12'd471  : out_data_ref <= 8'hdd;
      12'd472  : out_data_ref <= 8'hcc;
      12'd473  : out_data_ref <= 8'h52;
      12'd474  : out_data_ref <= 8'hbc;
      12'd475  : out_data_ref <= 8'h45;
      12'd476  : out_data_ref <= 8'hd4;
      12'd477  : out_data_ref <= 8'h81;
      12'd478  : out_data_ref <= 8'hcd;
      12'd479  : out_data_ref <= 8'hcf;
      12'd480  : out_data_ref <= 8'h74;
      12'd481  : out_data_ref <= 8'h47;
      12'd482  : out_data_ref <= 8'h3a;
      12'd483  : out_data_ref <= 8'h4f;
      12'd484  : out_data_ref <= 8'he3;
      12'd485  : out_data_ref <= 8'h09;
      12'd486  : out_data_ref <= 8'he4;
      12'd487  : out_data_ref <= 8'h41;
      12'd488  : out_data_ref <= 8'hb8;
      12'd489  : out_data_ref <= 8'h98;
      12'd490  : out_data_ref <= 8'h41;
      12'd491  : out_data_ref <= 8'hee;
      12'd492  : out_data_ref <= 8'h43;
      12'd493  : out_data_ref <= 8'h27;
      12'd494  : out_data_ref <= 8'hd1;
      12'd495  : out_data_ref <= 8'h22;
      12'd496  : out_data_ref <= 8'h16;
      12'd497  : out_data_ref <= 8'hd4;
      12'd498  : out_data_ref <= 8'h52;
      12'd499  : out_data_ref <= 8'hc1;
      12'd500  : out_data_ref <= 8'hda;
      12'd501  : out_data_ref <= 8'hcb;
      12'd502  : out_data_ref <= 8'hcb;
      12'd503  : out_data_ref <= 8'h6a;
      12'd504  : out_data_ref <= 8'h19;
      12'd505  : out_data_ref <= 8'h31;
      12'd506  : out_data_ref <= 8'h2c;
      12'd507  : out_data_ref <= 8'h3a;
      12'd508  : out_data_ref <= 8'ha7;
      12'd509  : out_data_ref <= 8'hdf;
      12'd510  : out_data_ref <= 8'h9e;
      12'd511  : out_data_ref <= 8'h52;
      12'd512  : out_data_ref <= 8'h0e;
      12'd513  : out_data_ref <= 8'h3b;
      12'd514  : out_data_ref <= 8'h37;
      12'd515  : out_data_ref <= 8'h61;
      12'd516  : out_data_ref <= 8'h92;
      12'd517  : out_data_ref <= 8'h33;
      12'd518  : out_data_ref <= 8'h33;
      12'd519  : out_data_ref <= 8'h18;
      12'd520  : out_data_ref <= 8'h12;
      12'd521  : out_data_ref <= 8'h26;
      12'd522  : out_data_ref <= 8'hf7;
      12'd523  : out_data_ref <= 8'h51;
      12'd524  : out_data_ref <= 8'he7;
      12'd525  : out_data_ref <= 8'h6c;
      12'd526  : out_data_ref <= 8'hb0;
      12'd527  : out_data_ref <= 8'h16;
      12'd528  : out_data_ref <= 8'hb6;
      12'd529  : out_data_ref <= 8'h5f;
      12'd530  : out_data_ref <= 8'h47;
      12'd531  : out_data_ref <= 8'h7f;
      12'd532  : out_data_ref <= 8'hbe;
      12'd533  : out_data_ref <= 8'h8f;
      12'd534  : out_data_ref <= 8'h6e;
      12'd535  : out_data_ref <= 8'hbc;
      12'd536  : out_data_ref <= 8'hb3;
      12'd537  : out_data_ref <= 8'h3d;
      12'd538  : out_data_ref <= 8'h36;
      12'd539  : out_data_ref <= 8'hf3;
      12'd540  : out_data_ref <= 8'ha5;
      12'd541  : out_data_ref <= 8'h6b;
      12'd542  : out_data_ref <= 8'h06;
      12'd543  : out_data_ref <= 8'hc9;
      12'd544  : out_data_ref <= 8'ha2;
      12'd545  : out_data_ref <= 8'he0;
      12'd546  : out_data_ref <= 8'h1c;
      12'd547  : out_data_ref <= 8'h3a;
      12'd548  : out_data_ref <= 8'h8a;
      12'd549  : out_data_ref <= 8'h8d;
      12'd550  : out_data_ref <= 8'h9c;
      12'd551  : out_data_ref <= 8'hb4;
      12'd552  : out_data_ref <= 8'h72;
      12'd553  : out_data_ref <= 8'h99;
      12'd554  : out_data_ref <= 8'hf2;
      12'd555  : out_data_ref <= 8'h18;
      12'd556  : out_data_ref <= 8'h3d;
      12'd557  : out_data_ref <= 8'ha8;
      12'd558  : out_data_ref <= 8'h17;
      12'd559  : out_data_ref <= 8'had;
      12'd560  : out_data_ref <= 8'h4c;
      12'd561  : out_data_ref <= 8'hfa;
      12'd562  : out_data_ref <= 8'h86;
      12'd563  : out_data_ref <= 8'h17;
      12'd564  : out_data_ref <= 8'h6e;
      12'd565  : out_data_ref <= 8'ha3;
      12'd566  : out_data_ref <= 8'hf7;
      12'd567  : out_data_ref <= 8'he3;
      12'd568  : out_data_ref <= 8'he1;
      12'd569  : out_data_ref <= 8'h1a;
      12'd570  : out_data_ref <= 8'he4;
      12'd571  : out_data_ref <= 8'h56;
      12'd572  : out_data_ref <= 8'hb1;
      12'd573  : out_data_ref <= 8'he4;
      12'd574  : out_data_ref <= 8'h11;
      12'd575  : out_data_ref <= 8'h24;
      12'd576  : out_data_ref <= 8'h71;
      12'd577  : out_data_ref <= 8'hb1;
      12'd578  : out_data_ref <= 8'ha1;
      12'd579  : out_data_ref <= 8'h55;
      12'd580  : out_data_ref <= 8'hc4;
      12'd581  : out_data_ref <= 8'h49;
      12'd582  : out_data_ref <= 8'h23;
      12'd583  : out_data_ref <= 8'h22;
      12'd584  : out_data_ref <= 8'h43;
      12'd585  : out_data_ref <= 8'h74;
      12'd586  : out_data_ref <= 8'hed;
      12'd587  : out_data_ref <= 8'h50;
      12'd588  : out_data_ref <= 8'h28;
      12'd589  : out_data_ref <= 8'h89;
      12'd590  : out_data_ref <= 8'h1e;
      12'd591  : out_data_ref <= 8'h1a;
      12'd592  : out_data_ref <= 8'h8d;
      12'd593  : out_data_ref <= 8'h2b;
      12'd594  : out_data_ref <= 8'hc6;
      12'd595  : out_data_ref <= 8'hec;
      12'd596  : out_data_ref <= 8'ha6;
      12'd597  : out_data_ref <= 8'h05;
      12'd598  : out_data_ref <= 8'ha8;
      12'd599  : out_data_ref <= 8'h17;
      12'd600  : out_data_ref <= 8'he1;
      12'd601  : out_data_ref <= 8'h6e;
      12'd602  : out_data_ref <= 8'hd2;
      12'd603  : out_data_ref <= 8'heb;
      12'd604  : out_data_ref <= 8'h12;
      12'd605  : out_data_ref <= 8'hcb;
      12'd606  : out_data_ref <= 8'h67;
      12'd607  : out_data_ref <= 8'hd1;
      12'd608  : out_data_ref <= 8'h71;
      12'd609  : out_data_ref <= 8'h1f;
      12'd610  : out_data_ref <= 8'hd8;
      12'd611  : out_data_ref <= 8'h6d;
      12'd612  : out_data_ref <= 8'h59;
      12'd613  : out_data_ref <= 8'h0b;
      12'd614  : out_data_ref <= 8'h2a;
      12'd615  : out_data_ref <= 8'h4d;
      12'd616  : out_data_ref <= 8'h56;
      12'd617  : out_data_ref <= 8'hd7;
      12'd618  : out_data_ref <= 8'h70;
      12'd619  : out_data_ref <= 8'hc4;
      12'd620  : out_data_ref <= 8'h4c;
      12'd621  : out_data_ref <= 8'he5;
      12'd622  : out_data_ref <= 8'hae;
      12'd623  : out_data_ref <= 8'hb3;
      12'd624  : out_data_ref <= 8'h7a;
      12'd625  : out_data_ref <= 8'hcd;
      12'd626  : out_data_ref <= 8'hd9;
      12'd627  : out_data_ref <= 8'hc4;
      12'd628  : out_data_ref <= 8'h39;
      12'd629  : out_data_ref <= 8'h17;
      12'd630  : out_data_ref <= 8'h64;
      12'd631  : out_data_ref <= 8'hbd;
      12'd632  : out_data_ref <= 8'h5d;
      12'd633  : out_data_ref <= 8'ha3;
      12'd634  : out_data_ref <= 8'h6c;
      12'd635  : out_data_ref <= 8'h2a;
      12'd636  : out_data_ref <= 8'h07;
      12'd637  : out_data_ref <= 8'hf4;
      12'd638  : out_data_ref <= 8'hcf;
      12'd639  : out_data_ref <= 8'he4;
      12'd640  : out_data_ref <= 8'h8c;
      12'd641  : out_data_ref <= 8'hae;
      12'd642  : out_data_ref <= 8'h24;
      12'd643  : out_data_ref <= 8'h41;
      12'd644  : out_data_ref <= 8'h4b;
      12'd645  : out_data_ref <= 8'h87;
      12'd646  : out_data_ref <= 8'he7;
      12'd647  : out_data_ref <= 8'h8d;
      12'd648  : out_data_ref <= 8'hb8;
      12'd649  : out_data_ref <= 8'h37;
      12'd650  : out_data_ref <= 8'h73;
      12'd651  : out_data_ref <= 8'h0e;
      12'd652  : out_data_ref <= 8'ha6;
      12'd653  : out_data_ref <= 8'h17;
      12'd654  : out_data_ref <= 8'hd2;
      12'd655  : out_data_ref <= 8'hb9;
      12'd656  : out_data_ref <= 8'hc8;
      12'd657  : out_data_ref <= 8'h28;
      12'd658  : out_data_ref <= 8'hc9;
      12'd659  : out_data_ref <= 8'h97;
      12'd660  : out_data_ref <= 8'h13;
      12'd661  : out_data_ref <= 8'h64;
      12'd662  : out_data_ref <= 8'h0f;
      12'd663  : out_data_ref <= 8'h10;
      12'd664  : out_data_ref <= 8'hae;
      12'd665  : out_data_ref <= 8'hf6;
      12'd666  : out_data_ref <= 8'hdf;
      12'd667  : out_data_ref <= 8'h80;
      12'd668  : out_data_ref <= 8'h37;
      12'd669  : out_data_ref <= 8'hc1;
      12'd670  : out_data_ref <= 8'h51;
      12'd671  : out_data_ref <= 8'hee;
      12'd672  : out_data_ref <= 8'h55;
      12'd673  : out_data_ref <= 8'h02;
      12'd674  : out_data_ref <= 8'hb5;
      12'd675  : out_data_ref <= 8'h27;
      12'd676  : out_data_ref <= 8'h29;
      12'd677  : out_data_ref <= 8'hc1;
      12'd678  : out_data_ref <= 8'hee;
      12'd679  : out_data_ref <= 8'hf4;
      12'd680  : out_data_ref <= 8'h60;
      12'd681  : out_data_ref <= 8'hde;
      12'd682  : out_data_ref <= 8'hca;
      12'd683  : out_data_ref <= 8'hed;
      12'd684  : out_data_ref <= 8'h3c;
      12'd685  : out_data_ref <= 8'hf4;
      12'd686  : out_data_ref <= 8'h71;
      12'd687  : out_data_ref <= 8'h76;
      12'd688  : out_data_ref <= 8'hd7;
      12'd689  : out_data_ref <= 8'h68;
      12'd690  : out_data_ref <= 8'hb4;
      12'd691  : out_data_ref <= 8'hf1;
      12'd692  : out_data_ref <= 8'hfc;
      12'd693  : out_data_ref <= 8'h47;
      12'd694  : out_data_ref <= 8'h5a;
      12'd695  : out_data_ref <= 8'h0f;
      12'd696  : out_data_ref <= 8'h8a;
      12'd697  : out_data_ref <= 8'h10;
      12'd698  : out_data_ref <= 8'h1d;
      12'd699  : out_data_ref <= 8'hcd;
      12'd700  : out_data_ref <= 8'hef;
      12'd701  : out_data_ref <= 8'he1;
      12'd702  : out_data_ref <= 8'h36;
      12'd703  : out_data_ref <= 8'h69;
      12'd704  : out_data_ref <= 8'h53;
      12'd705  : out_data_ref <= 8'h9d;
      12'd706  : out_data_ref <= 8'h91;
      12'd707  : out_data_ref <= 8'he8;
      12'd708  : out_data_ref <= 8'hda;
      12'd709  : out_data_ref <= 8'h0d;
      12'd710  : out_data_ref <= 8'h7e;
      12'd711  : out_data_ref <= 8'he9;
      12'd712  : out_data_ref <= 8'h6c;
      12'd713  : out_data_ref <= 8'hf3;
      12'd714  : out_data_ref <= 8'hc4;
      12'd715  : out_data_ref <= 8'hc5;
      12'd716  : out_data_ref <= 8'hb0;
      12'd717  : out_data_ref <= 8'h31;
      12'd718  : out_data_ref <= 8'h86;
      12'd719  : out_data_ref <= 8'h3a;
      12'd720  : out_data_ref <= 8'hc3;
      12'd721  : out_data_ref <= 8'hd1;
      12'd722  : out_data_ref <= 8'hae;
      12'd723  : out_data_ref <= 8'h7c;
      12'd724  : out_data_ref <= 8'hb0;
      12'd725  : out_data_ref <= 8'h7b;
      12'd726  : out_data_ref <= 8'h81;
      12'd727  : out_data_ref <= 8'h3f;
      12'd728  : out_data_ref <= 8'h7f;
      12'd729  : out_data_ref <= 8'h1b;
      12'd730  : out_data_ref <= 8'h2c;
      12'd731  : out_data_ref <= 8'hb3;
      12'd732  : out_data_ref <= 8'h4f;
      12'd733  : out_data_ref <= 8'he4;
      12'd734  : out_data_ref <= 8'h17;
      12'd735  : out_data_ref <= 8'h92;
      12'd736  : out_data_ref <= 8'hf1;
      12'd737  : out_data_ref <= 8'h19;
      12'd738  : out_data_ref <= 8'hf8;
      12'd739  : out_data_ref <= 8'hbf;
      12'd740  : out_data_ref <= 8'h11;
      12'd741  : out_data_ref <= 8'h32;
      12'd742  : out_data_ref <= 8'hd8;
      12'd743  : out_data_ref <= 8'hbe;
      12'd744  : out_data_ref <= 8'hee;
      12'd745  : out_data_ref <= 8'h77;
      12'd746  : out_data_ref <= 8'h54;
      12'd747  : out_data_ref <= 8'h41;
      12'd748  : out_data_ref <= 8'hfd;
      12'd749  : out_data_ref <= 8'h0f;
      12'd750  : out_data_ref <= 8'h95;
      12'd751  : out_data_ref <= 8'h42;
      12'd752  : out_data_ref <= 8'h16;
      12'd753  : out_data_ref <= 8'h60;
      12'd754  : out_data_ref <= 8'h5a;
      12'd755  : out_data_ref <= 8'hb8;
      12'd756  : out_data_ref <= 8'h52;
      12'd757  : out_data_ref <= 8'h79;
      12'd758  : out_data_ref <= 8'h7d;
      12'd759  : out_data_ref <= 8'h09;
      12'd760  : out_data_ref <= 8'h02;
      12'd761  : out_data_ref <= 8'hce;
      12'd762  : out_data_ref <= 8'h9b;
      12'd763  : out_data_ref <= 8'h30;
      12'd764  : out_data_ref <= 8'h4c;
      12'd765  : out_data_ref <= 8'h7d;
      12'd766  : out_data_ref <= 8'h34;
      12'd767  : out_data_ref <= 8'h38;
      12'd768  : out_data_ref <= 8'h82;
      12'd769  : out_data_ref <= 8'h0c;
      12'd770  : out_data_ref <= 8'h48;
      12'd771  : out_data_ref <= 8'h5d;
      12'd772  : out_data_ref <= 8'h2c;
      12'd773  : out_data_ref <= 8'h2e;
      12'd774  : out_data_ref <= 8'hbb;
      12'd775  : out_data_ref <= 8'h0a;
      12'd776  : out_data_ref <= 8'hda;
      12'd777  : out_data_ref <= 8'he3;
      12'd778  : out_data_ref <= 8'he0;
      12'd779  : out_data_ref <= 8'h31;
      12'd780  : out_data_ref <= 8'h7e;
      12'd781  : out_data_ref <= 8'h55;
      12'd782  : out_data_ref <= 8'h68;
      12'd783  : out_data_ref <= 8'h83;
      12'd784  : out_data_ref <= 8'h13;
      12'd785  : out_data_ref <= 8'hf2;
      12'd786  : out_data_ref <= 8'hd1;
      12'd787  : out_data_ref <= 8'h18;
      12'd788  : out_data_ref <= 8'h4e;
      12'd789  : out_data_ref <= 8'he1;
      12'd790  : out_data_ref <= 8'hd8;
      12'd791  : out_data_ref <= 8'h6e;
      12'd792  : out_data_ref <= 8'h81;
      12'd793  : out_data_ref <= 8'had;
      12'd794  : out_data_ref <= 8'heb;
      12'd795  : out_data_ref <= 8'h36;
      12'd796  : out_data_ref <= 8'h55;
      12'd797  : out_data_ref <= 8'h5d;
      12'd798  : out_data_ref <= 8'h7e;
      12'd799  : out_data_ref <= 8'h22;
      12'd800  : out_data_ref <= 8'h54;
      12'd801  : out_data_ref <= 8'h0b;
      12'd802  : out_data_ref <= 8'h38;
      12'd803  : out_data_ref <= 8'h1a;
      12'd804  : out_data_ref <= 8'h03;
      12'd805  : out_data_ref <= 8'h87;
      12'd806  : out_data_ref <= 8'h2b;
      12'd807  : out_data_ref <= 8'h66;
      12'd808  : out_data_ref <= 8'hd7;
      12'd809  : out_data_ref <= 8'hb8;
      12'd810  : out_data_ref <= 8'hae;
      12'd811  : out_data_ref <= 8'hf9;
      12'd812  : out_data_ref <= 8'h75;
      12'd813  : out_data_ref <= 8'h81;
      12'd814  : out_data_ref <= 8'h94;
      12'd815  : out_data_ref <= 8'h3f;
      12'd816  : out_data_ref <= 8'h67;
      12'd817  : out_data_ref <= 8'hdf;
      12'd818  : out_data_ref <= 8'he4;
      12'd819  : out_data_ref <= 8'h27;
      12'd820  : out_data_ref <= 8'hea;
      12'd821  : out_data_ref <= 8'h64;
      12'd822  : out_data_ref <= 8'h24;
      12'd823  : out_data_ref <= 8'h67;
      12'd824  : out_data_ref <= 8'h25;
      12'd825  : out_data_ref <= 8'h45;
      12'd826  : out_data_ref <= 8'ha6;
      12'd827  : out_data_ref <= 8'hc9;
      12'd828  : out_data_ref <= 8'h5d;
      12'd829  : out_data_ref <= 8'hd0;
      12'd830  : out_data_ref <= 8'h32;
      12'd831  : out_data_ref <= 8'h0d;
      12'd832  : out_data_ref <= 8'h16;
      12'd833  : out_data_ref <= 8'h13;
      12'd834  : out_data_ref <= 8'hd0;
      12'd835  : out_data_ref <= 8'h65;
      12'd836  : out_data_ref <= 8'h82;
      12'd837  : out_data_ref <= 8'h2b;
      12'd838  : out_data_ref <= 8'h8f;
      12'd839  : out_data_ref <= 8'h15;
      12'd840  : out_data_ref <= 8'h6f;
      12'd841  : out_data_ref <= 8'h67;
      12'd842  : out_data_ref <= 8'h1f;
      12'd843  : out_data_ref <= 8'h78;
      12'd844  : out_data_ref <= 8'hfe;
      12'd845  : out_data_ref <= 8'h75;
      12'd846  : out_data_ref <= 8'hf5;
      12'd847  : out_data_ref <= 8'h60;
      12'd848  : out_data_ref <= 8'hdd;
      12'd849  : out_data_ref <= 8'he7;
      12'd850  : out_data_ref <= 8'h67;
      12'd851  : out_data_ref <= 8'h4d;
      12'd852  : out_data_ref <= 8'hc9;
      12'd853  : out_data_ref <= 8'hc1;
      12'd854  : out_data_ref <= 8'h53;
      12'd855  : out_data_ref <= 8'h61;
      12'd856  : out_data_ref <= 8'h79;
      12'd857  : out_data_ref <= 8'hda;
      12'd858  : out_data_ref <= 8'h1a;
      12'd859  : out_data_ref <= 8'hbe;
      12'd860  : out_data_ref <= 8'hfb;
      12'd861  : out_data_ref <= 8'h30;
      12'd862  : out_data_ref <= 8'haa;
      12'd863  : out_data_ref <= 8'h54;
      12'd864  : out_data_ref <= 8'h56;
      12'd865  : out_data_ref <= 8'h1c;
      12'd866  : out_data_ref <= 8'hf2;
      12'd867  : out_data_ref <= 8'hfa;
      12'd868  : out_data_ref <= 8'hdb;
      12'd869  : out_data_ref <= 8'h39;
      12'd870  : out_data_ref <= 8'h28;
      12'd871  : out_data_ref <= 8'h2f;
      12'd872  : out_data_ref <= 8'h94;
      12'd873  : out_data_ref <= 8'hae;
      12'd874  : out_data_ref <= 8'ha3;
      12'd875  : out_data_ref <= 8'h3f;
      12'd876  : out_data_ref <= 8'h19;
      12'd877  : out_data_ref <= 8'h41;
      12'd878  : out_data_ref <= 8'h96;
      12'd879  : out_data_ref <= 8'hd2;
      12'd880  : out_data_ref <= 8'h6d;
      12'd881  : out_data_ref <= 8'hd6;
      12'd882  : out_data_ref <= 8'h5c;
      12'd883  : out_data_ref <= 8'hd6;
      12'd884  : out_data_ref <= 8'h5d;
      12'd885  : out_data_ref <= 8'hcd;
      12'd886  : out_data_ref <= 8'h70;
      12'd887  : out_data_ref <= 8'ha4;
      12'd888  : out_data_ref <= 8'h08;
      12'd889  : out_data_ref <= 8'h6f;
      12'd890  : out_data_ref <= 8'h9e;
      12'd891  : out_data_ref <= 8'h35;
      12'd892  : out_data_ref <= 8'h58;
      12'd893  : out_data_ref <= 8'h09;
      12'd894  : out_data_ref <= 8'hdc;
      12'd895  : out_data_ref <= 8'h27;
      12'd896  : out_data_ref <= 8'h01;
      12'd897  : out_data_ref <= 8'h9c;
      12'd898  : out_data_ref <= 8'he6;
      12'd899  : out_data_ref <= 8'h91;
      12'd900  : out_data_ref <= 8'hd5;
      12'd901  : out_data_ref <= 8'h02;
      12'd902  : out_data_ref <= 8'he6;
      12'd903  : out_data_ref <= 8'h7f;
      12'd904  : out_data_ref <= 8'h55;
      12'd905  : out_data_ref <= 8'h3e;
      12'd906  : out_data_ref <= 8'h25;
      12'd907  : out_data_ref <= 8'hb9;
      12'd908  : out_data_ref <= 8'h69;
      12'd909  : out_data_ref <= 8'h54;
      12'd910  : out_data_ref <= 8'h51;
      12'd911  : out_data_ref <= 8'hce;
      12'd912  : out_data_ref <= 8'hbb;
      12'd913  : out_data_ref <= 8'he6;
      12'd914  : out_data_ref <= 8'hdb;
      12'd915  : out_data_ref <= 8'h28;
      12'd916  : out_data_ref <= 8'h53;
      12'd917  : out_data_ref <= 8'h8d;
      12'd918  : out_data_ref <= 8'h34;
      12'd919  : out_data_ref <= 8'hcd;
      12'd920  : out_data_ref <= 8'h08;
      12'd921  : out_data_ref <= 8'h4e;
      12'd922  : out_data_ref <= 8'h41;
      12'd923  : out_data_ref <= 8'h5a;
      12'd924  : out_data_ref <= 8'h74;
      12'd925  : out_data_ref <= 8'h65;
      12'd926  : out_data_ref <= 8'h12;
      12'd927  : out_data_ref <= 8'h36;
      12'd928  : out_data_ref <= 8'h08;
      12'd929  : out_data_ref <= 8'h8a;
      12'd930  : out_data_ref <= 8'h10;
      12'd931  : out_data_ref <= 8'hbd;
      12'd932  : out_data_ref <= 8'h00;
      12'd933  : out_data_ref <= 8'hbe;
      12'd934  : out_data_ref <= 8'h53;
      12'd935  : out_data_ref <= 8'h41;
      12'd936  : out_data_ref <= 8'h3a;
      12'd937  : out_data_ref <= 8'hd1;
      12'd938  : out_data_ref <= 8'h24;
      12'd939  : out_data_ref <= 8'h9a;
      12'd940  : out_data_ref <= 8'hab;
      12'd941  : out_data_ref <= 8'hb2;
      12'd942  : out_data_ref <= 8'h2b;
      12'd943  : out_data_ref <= 8'hd3;
      12'd944  : out_data_ref <= 8'h99;
      12'd945  : out_data_ref <= 8'h7e;
      12'd946  : out_data_ref <= 8'h10;
      12'd947  : out_data_ref <= 8'h3b;
      12'd948  : out_data_ref <= 8'hea;
      12'd949  : out_data_ref <= 8'h45;
      12'd950  : out_data_ref <= 8'h93;
      12'd951  : out_data_ref <= 8'h82;
      12'd952  : out_data_ref <= 8'h06;
      12'd953  : out_data_ref <= 8'hcf;
      12'd954  : out_data_ref <= 8'h68;
      12'd955  : out_data_ref <= 8'h51;
      12'd956  : out_data_ref <= 8'h4b;
      12'd957  : out_data_ref <= 8'h58;
      12'd958  : out_data_ref <= 8'h24;
      12'd959  : out_data_ref <= 8'h27;
      12'd960  : out_data_ref <= 8'hcf;
      12'd961  : out_data_ref <= 8'h00;
      12'd962  : out_data_ref <= 8'h98;
      12'd963  : out_data_ref <= 8'h57;
      12'd964  : out_data_ref <= 8'hab;
      12'd965  : out_data_ref <= 8'h20;
      12'd966  : out_data_ref <= 8'h8f;
      12'd967  : out_data_ref <= 8'h59;
      12'd968  : out_data_ref <= 8'he2;
      12'd969  : out_data_ref <= 8'h23;
      12'd970  : out_data_ref <= 8'hf8;
      12'd971  : out_data_ref <= 8'hfc;
      12'd972  : out_data_ref <= 8'h02;
      12'd973  : out_data_ref <= 8'he4;
      12'd974  : out_data_ref <= 8'h16;
      12'd975  : out_data_ref <= 8'h62;
      12'd976  : out_data_ref <= 8'hc5;
      12'd977  : out_data_ref <= 8'h05;
      12'd978  : out_data_ref <= 8'ha2;
      12'd979  : out_data_ref <= 8'h97;
      12'd980  : out_data_ref <= 8'h32;
      12'd981  : out_data_ref <= 8'ha8;
      12'd982  : out_data_ref <= 8'h42;
      12'd983  : out_data_ref <= 8'h18;
      12'd984  : out_data_ref <= 8'h70;
      12'd985  : out_data_ref <= 8'h56;
      12'd986  : out_data_ref <= 8'h69;
      12'd987  : out_data_ref <= 8'hf9;
      12'd988  : out_data_ref <= 8'h09;
      12'd989  : out_data_ref <= 8'hfc;
      12'd990  : out_data_ref <= 8'hb1;
      12'd991  : out_data_ref <= 8'h27;
      12'd992  : out_data_ref <= 8'hb4;
      12'd993  : out_data_ref <= 8'h0b;
      12'd994  : out_data_ref <= 8'h82;
      12'd995  : out_data_ref <= 8'h74;
      12'd996  : out_data_ref <= 8'h7b;
      12'd997  : out_data_ref <= 8'h08;
      12'd998  : out_data_ref <= 8'h10;
      12'd999  : out_data_ref <= 8'h21;
      12'd1000 : out_data_ref <= 8'h53;
      12'd1001 : out_data_ref <= 8'h71;
      12'd1002 : out_data_ref <= 8'h0b;
      12'd1003 : out_data_ref <= 8'h8c;
      12'd1004 : out_data_ref <= 8'hc9;
      12'd1005 : out_data_ref <= 8'h5a;
      12'd1006 : out_data_ref <= 8'h3b;
      12'd1007 : out_data_ref <= 8'h7a;
      12'd1008 : out_data_ref <= 8'hbc;
      12'd1009 : out_data_ref <= 8'h0d;
      12'd1010 : out_data_ref <= 8'hd4;
      12'd1011 : out_data_ref <= 8'h01;
      12'd1012 : out_data_ref <= 8'h15;
      12'd1013 : out_data_ref <= 8'h83;
      12'd1014 : out_data_ref <= 8'hed;
      12'd1015 : out_data_ref <= 8'ha3;
      12'd1016 : out_data_ref <= 8'h59;
      12'd1017 : out_data_ref <= 8'h82;
      12'd1018 : out_data_ref <= 8'hfc;
      12'd1019 : out_data_ref <= 8'hf2;
      12'd1020 : out_data_ref <= 8'h0d;
      12'd1021 : out_data_ref <= 8'h95;
      12'd1022 : out_data_ref <= 8'he5;
      12'd1023 : out_data_ref <= 8'h87;
      12'd1024 : out_data_ref <= 8'h3c;
      12'd1025 : out_data_ref <= 8'h7a;
      12'd1026 : out_data_ref <= 8'h97;
      12'd1027 : out_data_ref <= 8'h63;
      12'd1028 : out_data_ref <= 8'hd9;
      12'd1029 : out_data_ref <= 8'hd0;
      12'd1030 : out_data_ref <= 8'hf9;
      12'd1031 : out_data_ref <= 8'h10;
      12'd1032 : out_data_ref <= 8'h88;
      12'd1033 : out_data_ref <= 8'hbb;
      12'd1034 : out_data_ref <= 8'hdf;
      12'd1035 : out_data_ref <= 8'h07;
      12'd1036 : out_data_ref <= 8'h1f;
      12'd1037 : out_data_ref <= 8'h10;
      12'd1038 : out_data_ref <= 8'h8d;
      12'd1039 : out_data_ref <= 8'h89;
      12'd1040 : out_data_ref <= 8'he6;
      12'd1041 : out_data_ref <= 8'h6d;
      12'd1042 : out_data_ref <= 8'h20;
      12'd1043 : out_data_ref <= 8'hbc;
      12'd1044 : out_data_ref <= 8'hef;
      12'd1045 : out_data_ref <= 8'hca;
      12'd1046 : out_data_ref <= 8'h8b;
      12'd1047 : out_data_ref <= 8'hd6;
      12'd1048 : out_data_ref <= 8'h61;
      12'd1049 : out_data_ref <= 8'h3d;
      12'd1050 : out_data_ref <= 8'hfa;
      12'd1051 : out_data_ref <= 8'h38;
      12'd1052 : out_data_ref <= 8'h9d;
      12'd1053 : out_data_ref <= 8'hbe;
      12'd1054 : out_data_ref <= 8'hed;
      12'd1055 : out_data_ref <= 8'hb2;
      12'd1056 : out_data_ref <= 8'h6d;
      12'd1057 : out_data_ref <= 8'h23;
      12'd1058 : out_data_ref <= 8'hbf;
      12'd1059 : out_data_ref <= 8'h50;
      12'd1060 : out_data_ref <= 8'h00;
      12'd1061 : out_data_ref <= 8'h06;
      12'd1062 : out_data_ref <= 8'h8b;
      12'd1063 : out_data_ref <= 8'hfb;
      12'd1064 : out_data_ref <= 8'h76;
      12'd1065 : out_data_ref <= 8'hd2;
      12'd1066 : out_data_ref <= 8'h9e;
      12'd1067 : out_data_ref <= 8'hb8;
      12'd1068 : out_data_ref <= 8'h65;
      12'd1069 : out_data_ref <= 8'hf6;
      12'd1070 : out_data_ref <= 8'h3d;
      12'd1071 : out_data_ref <= 8'h9a;
      12'd1072 : out_data_ref <= 8'h45;
      12'd1073 : out_data_ref <= 8'hb1;
      12'd1074 : out_data_ref <= 8'hd4;
      12'd1075 : out_data_ref <= 8'hd8;
      12'd1076 : out_data_ref <= 8'h47;
      12'd1077 : out_data_ref <= 8'hba;
      12'd1078 : out_data_ref <= 8'h9d;
      12'd1079 : out_data_ref <= 8'h71;
      12'd1080 : out_data_ref <= 8'h68;
      12'd1081 : out_data_ref <= 8'hd0;
      12'd1082 : out_data_ref <= 8'h89;
      12'd1083 : out_data_ref <= 8'h3d;
      12'd1084 : out_data_ref <= 8'h13;
      12'd1085 : out_data_ref <= 8'h42;
      12'd1086 : out_data_ref <= 8'h6c;
      12'd1087 : out_data_ref <= 8'hd2;
      12'd1088 : out_data_ref <= 8'h8d;
      12'd1089 : out_data_ref <= 8'h3b;
      12'd1090 : out_data_ref <= 8'hb7;
      12'd1091 : out_data_ref <= 8'h4f;
      12'd1092 : out_data_ref <= 8'h21;
      12'd1093 : out_data_ref <= 8'hbe;
      12'd1094 : out_data_ref <= 8'hfe;
      12'd1095 : out_data_ref <= 8'h4a;
      12'd1096 : out_data_ref <= 8'h8b;
      12'd1097 : out_data_ref <= 8'he8;
      12'd1098 : out_data_ref <= 8'h6a;
      12'd1099 : out_data_ref <= 8'hc2;
      12'd1100 : out_data_ref <= 8'ha4;
      12'd1101 : out_data_ref <= 8'h55;
      12'd1102 : out_data_ref <= 8'hbd;
      12'd1103 : out_data_ref <= 8'hd7;
      12'd1104 : out_data_ref <= 8'h01;
      12'd1105 : out_data_ref <= 8'h6f;
      12'd1106 : out_data_ref <= 8'h38;
      12'd1107 : out_data_ref <= 8'hac;
      12'd1108 : out_data_ref <= 8'h0c;
      12'd1109 : out_data_ref <= 8'h62;
      12'd1110 : out_data_ref <= 8'hdb;
      12'd1111 : out_data_ref <= 8'h66;
      12'd1112 : out_data_ref <= 8'hc0;
      12'd1113 : out_data_ref <= 8'h25;
      12'd1114 : out_data_ref <= 8'hfd;
      12'd1115 : out_data_ref <= 8'h89;
      12'd1116 : out_data_ref <= 8'h04;
      12'd1117 : out_data_ref <= 8'hf0;
      12'd1118 : out_data_ref <= 8'h22;
      12'd1119 : out_data_ref <= 8'h7e;
      12'd1120 : out_data_ref <= 8'hf6;
      12'd1121 : out_data_ref <= 8'hbd;
      12'd1122 : out_data_ref <= 8'hd7;
      12'd1123 : out_data_ref <= 8'h06;
      12'd1124 : out_data_ref <= 8'h9a;
      12'd1125 : out_data_ref <= 8'h2c;
      12'd1126 : out_data_ref <= 8'h7d;
      12'd1127 : out_data_ref <= 8'h53;
      12'd1128 : out_data_ref <= 8'h5d;
      12'd1129 : out_data_ref <= 8'hd8;
      12'd1130 : out_data_ref <= 8'hd3;
      12'd1131 : out_data_ref <= 8'h55;
      12'd1132 : out_data_ref <= 8'h5f;
      12'd1133 : out_data_ref <= 8'h08;
      12'd1134 : out_data_ref <= 8'h7f;
      12'd1135 : out_data_ref <= 8'h7c;
      12'd1136 : out_data_ref <= 8'h4c;
      12'd1137 : out_data_ref <= 8'h54;
      12'd1138 : out_data_ref <= 8'h8a;
      12'd1139 : out_data_ref <= 8'h03;
      12'd1140 : out_data_ref <= 8'ha2;
      12'd1141 : out_data_ref <= 8'hae;
      12'd1142 : out_data_ref <= 8'ha1;
      12'd1143 : out_data_ref <= 8'h41;
      12'd1144 : out_data_ref <= 8'h85;
      12'd1145 : out_data_ref <= 8'ha4;
      12'd1146 : out_data_ref <= 8'h9d;
      12'd1147 : out_data_ref <= 8'h18;
      12'd1148 : out_data_ref <= 8'h22;
      12'd1149 : out_data_ref <= 8'hed;
      12'd1150 : out_data_ref <= 8'h29;
      12'd1151 : out_data_ref <= 8'h79;
      12'd1152 : out_data_ref <= 8'h26;
      12'd1153 : out_data_ref <= 8'h5a;
      12'd1154 : out_data_ref <= 8'he0;
      12'd1155 : out_data_ref <= 8'h9f;
      12'd1156 : out_data_ref <= 8'h79;
      12'd1157 : out_data_ref <= 8'ha4;
      12'd1158 : out_data_ref <= 8'h43;
      12'd1159 : out_data_ref <= 8'hd3;
      12'd1160 : out_data_ref <= 8'hd7;
      12'd1161 : out_data_ref <= 8'he8;
      12'd1162 : out_data_ref <= 8'h20;
      12'd1163 : out_data_ref <= 8'h4f;
      12'd1164 : out_data_ref <= 8'hea;
      12'd1165 : out_data_ref <= 8'hb4;
      12'd1166 : out_data_ref <= 8'he9;
      12'd1167 : out_data_ref <= 8'h2b;
      12'd1168 : out_data_ref <= 8'h29;
      12'd1169 : out_data_ref <= 8'he7;
      12'd1170 : out_data_ref <= 8'he4;
      12'd1171 : out_data_ref <= 8'hb7;
      12'd1172 : out_data_ref <= 8'hbf;
      12'd1173 : out_data_ref <= 8'h18;
      12'd1174 : out_data_ref <= 8'h6f;
      12'd1175 : out_data_ref <= 8'h02;
      12'd1176 : out_data_ref <= 8'h43;
      12'd1177 : out_data_ref <= 8'h20;
      12'd1178 : out_data_ref <= 8'h9b;
      12'd1179 : out_data_ref <= 8'h92;
      12'd1180 : out_data_ref <= 8'h8b;
      12'd1181 : out_data_ref <= 8'h82;
      12'd1182 : out_data_ref <= 8'h38;
      12'd1183 : out_data_ref <= 8'ha1;
      12'd1184 : out_data_ref <= 8'h5e;
      12'd1185 : out_data_ref <= 8'h50;
      12'd1186 : out_data_ref <= 8'he9;
      12'd1187 : out_data_ref <= 8'h6a;
      12'd1188 : out_data_ref <= 8'h8c;
      12'd1189 : out_data_ref <= 8'h53;
      12'd1190 : out_data_ref <= 8'h7a;
      12'd1191 : out_data_ref <= 8'h44;
      12'd1192 : out_data_ref <= 8'h8f;
      12'd1193 : out_data_ref <= 8'hf2;
      12'd1194 : out_data_ref <= 8'he0;
      12'd1195 : out_data_ref <= 8'h88;
      12'd1196 : out_data_ref <= 8'hf9;
      12'd1197 : out_data_ref <= 8'h9f;
      12'd1198 : out_data_ref <= 8'hcb;
      12'd1199 : out_data_ref <= 8'h59;
      12'd1200 : out_data_ref <= 8'h02;
      12'd1201 : out_data_ref <= 8'hc8;
      12'd1202 : out_data_ref <= 8'h3b;
      12'd1203 : out_data_ref <= 8'h77;
      12'd1204 : out_data_ref <= 8'h6c;
      12'd1205 : out_data_ref <= 8'h1d;
      12'd1206 : out_data_ref <= 8'h09;
      12'd1207 : out_data_ref <= 8'h9d;
      12'd1208 : out_data_ref <= 8'h05;
      12'd1209 : out_data_ref <= 8'h69;
      12'd1210 : out_data_ref <= 8'hdb;
      12'd1211 : out_data_ref <= 8'hbf;
      12'd1212 : out_data_ref <= 8'h30;
      12'd1213 : out_data_ref <= 8'h27;
      12'd1214 : out_data_ref <= 8'ha4;
      12'd1215 : out_data_ref <= 8'h83;
      12'd1216 : out_data_ref <= 8'h64;
      12'd1217 : out_data_ref <= 8'hee;
      12'd1218 : out_data_ref <= 8'hb5;
      12'd1219 : out_data_ref <= 8'h11;
      12'd1220 : out_data_ref <= 8'hd3;
      12'd1221 : out_data_ref <= 8'h68;
      12'd1222 : out_data_ref <= 8'h4d;
      12'd1223 : out_data_ref <= 8'hba;
      12'd1224 : out_data_ref <= 8'h43;
      12'd1225 : out_data_ref <= 8'h4a;
      12'd1226 : out_data_ref <= 8'h92;
      12'd1227 : out_data_ref <= 8'h56;
      12'd1228 : out_data_ref <= 8'h0b;
      12'd1229 : out_data_ref <= 8'h37;
      12'd1230 : out_data_ref <= 8'h60;
      12'd1231 : out_data_ref <= 8'h64;
      12'd1232 : out_data_ref <= 8'h47;
      12'd1233 : out_data_ref <= 8'h36;
      12'd1234 : out_data_ref <= 8'h4a;
      12'd1235 : out_data_ref <= 8'hfa;
      12'd1236 : out_data_ref <= 8'h71;
      12'd1237 : out_data_ref <= 8'h87;
      12'd1238 : out_data_ref <= 8'h97;
      12'd1239 : out_data_ref <= 8'h89;
      12'd1240 : out_data_ref <= 8'hef;
      12'd1241 : out_data_ref <= 8'h88;
      12'd1242 : out_data_ref <= 8'hb7;
      12'd1243 : out_data_ref <= 8'hb4;
      12'd1244 : out_data_ref <= 8'h1f;
      12'd1245 : out_data_ref <= 8'h44;
      12'd1246 : out_data_ref <= 8'hd5;
      12'd1247 : out_data_ref <= 8'he0;
      12'd1248 : out_data_ref <= 8'h23;
      12'd1249 : out_data_ref <= 8'h7c;
      12'd1250 : out_data_ref <= 8'h8b;
      12'd1251 : out_data_ref <= 8'h92;
      12'd1252 : out_data_ref <= 8'h6c;
      12'd1253 : out_data_ref <= 8'hbe;
      12'd1254 : out_data_ref <= 8'h73;
      12'd1255 : out_data_ref <= 8'h9e;
      12'd1256 : out_data_ref <= 8'hd1;
      12'd1257 : out_data_ref <= 8'h5a;
      12'd1258 : out_data_ref <= 8'h57;
      12'd1259 : out_data_ref <= 8'h4a;
      12'd1260 : out_data_ref <= 8'had;
      12'd1261 : out_data_ref <= 8'hc5;
      12'd1262 : out_data_ref <= 8'h14;
      12'd1263 : out_data_ref <= 8'h7a;
      12'd1264 : out_data_ref <= 8'haa;
      12'd1265 : out_data_ref <= 8'h96;
      12'd1266 : out_data_ref <= 8'hd6;
      12'd1267 : out_data_ref <= 8'h12;
      12'd1268 : out_data_ref <= 8'h88;
      12'd1269 : out_data_ref <= 8'h8e;
      12'd1270 : out_data_ref <= 8'hbf;
      12'd1271 : out_data_ref <= 8'h4d;
      12'd1272 : out_data_ref <= 8'hf1;
      12'd1273 : out_data_ref <= 8'h24;
      12'd1274 : out_data_ref <= 8'h37;
      12'd1275 : out_data_ref <= 8'hbc;
      12'd1276 : out_data_ref <= 8'h9e;
      12'd1277 : out_data_ref <= 8'hd3;
      12'd1278 : out_data_ref <= 8'h3f;
      12'd1279 : out_data_ref <= 8'hab;
      12'd1280 : out_data_ref <= 8'hca;
      12'd1281 : out_data_ref <= 8'hd1;
      12'd1282 : out_data_ref <= 8'h8b;
      12'd1283 : out_data_ref <= 8'h3e;
      12'd1284 : out_data_ref <= 8'h1a;
      12'd1285 : out_data_ref <= 8'h0e;
      12'd1286 : out_data_ref <= 8'hbd;
      12'd1287 : out_data_ref <= 8'hb2;
      12'd1288 : out_data_ref <= 8'h1a;
      12'd1289 : out_data_ref <= 8'hfc;
      12'd1290 : out_data_ref <= 8'ha6;
      12'd1291 : out_data_ref <= 8'hfb;
      12'd1292 : out_data_ref <= 8'hd2;
      12'd1293 : out_data_ref <= 8'h71;
      12'd1294 : out_data_ref <= 8'h0b;
      12'd1295 : out_data_ref <= 8'h83;
      12'd1296 : out_data_ref <= 8'ha5;
      12'd1297 : out_data_ref <= 8'h57;
      12'd1298 : out_data_ref <= 8'h2d;
      12'd1299 : out_data_ref <= 8'hc8;
      12'd1300 : out_data_ref <= 8'h6a;
      12'd1301 : out_data_ref <= 8'h72;
      12'd1302 : out_data_ref <= 8'hf8;
      12'd1303 : out_data_ref <= 8'hff;
      12'd1304 : out_data_ref <= 8'h9a;
      12'd1305 : out_data_ref <= 8'h11;
      12'd1306 : out_data_ref <= 8'h5d;
      12'd1307 : out_data_ref <= 8'h82;
      12'd1308 : out_data_ref <= 8'h60;
      12'd1309 : out_data_ref <= 8'hd7;
      12'd1310 : out_data_ref <= 8'h90;
      12'd1311 : out_data_ref <= 8'h0f;
      12'd1312 : out_data_ref <= 8'he1;
      12'd1313 : out_data_ref <= 8'hf5;
      12'd1314 : out_data_ref <= 8'he1;
      12'd1315 : out_data_ref <= 8'h5e;
      12'd1316 : out_data_ref <= 8'h80;
      12'd1317 : out_data_ref <= 8'h7a;
      12'd1318 : out_data_ref <= 8'h20;
      12'd1319 : out_data_ref <= 8'h61;
      12'd1320 : out_data_ref <= 8'h8e;
      12'd1321 : out_data_ref <= 8'h0a;
      12'd1322 : out_data_ref <= 8'h75;
      12'd1323 : out_data_ref <= 8'he3;
      12'd1324 : out_data_ref <= 8'hfa;
      12'd1325 : out_data_ref <= 8'h5d;
      12'd1326 : out_data_ref <= 8'h4f;
      12'd1327 : out_data_ref <= 8'ha5;
      12'd1328 : out_data_ref <= 8'h97;
      12'd1329 : out_data_ref <= 8'h12;
      12'd1330 : out_data_ref <= 8'h89;
      12'd1331 : out_data_ref <= 8'h01;
      12'd1332 : out_data_ref <= 8'h24;
      12'd1333 : out_data_ref <= 8'h31;
      12'd1334 : out_data_ref <= 8'hc8;
      12'd1335 : out_data_ref <= 8'ha0;
      12'd1336 : out_data_ref <= 8'h35;
      12'd1337 : out_data_ref <= 8'hb5;
      12'd1338 : out_data_ref <= 8'hb2;
      12'd1339 : out_data_ref <= 8'hd7;
      12'd1340 : out_data_ref <= 8'hca;
      12'd1341 : out_data_ref <= 8'h0c;
      12'd1342 : out_data_ref <= 8'hf0;
      12'd1343 : out_data_ref <= 8'h46;
      12'd1344 : out_data_ref <= 8'hce;
      12'd1345 : out_data_ref <= 8'h79;
      12'd1346 : out_data_ref <= 8'h3a;
      12'd1347 : out_data_ref <= 8'ha4;
      12'd1348 : out_data_ref <= 8'h19;
      12'd1349 : out_data_ref <= 8'ha6;
      12'd1350 : out_data_ref <= 8'hb5;
      12'd1351 : out_data_ref <= 8'h8e;
      12'd1352 : out_data_ref <= 8'h4c;
      12'd1353 : out_data_ref <= 8'h77;
      12'd1354 : out_data_ref <= 8'hee;
      12'd1355 : out_data_ref <= 8'h5b;
      12'd1356 : out_data_ref <= 8'h2f;
      12'd1357 : out_data_ref <= 8'hf5;
      12'd1358 : out_data_ref <= 8'h48;
      12'd1359 : out_data_ref <= 8'h9c;
      12'd1360 : out_data_ref <= 8'hd0;
      12'd1361 : out_data_ref <= 8'hcd;
      12'd1362 : out_data_ref <= 8'hf5;
      12'd1363 : out_data_ref <= 8'h79;
      12'd1364 : out_data_ref <= 8'h07;
      12'd1365 : out_data_ref <= 8'h4f;
      12'd1366 : out_data_ref <= 8'h29;
      12'd1367 : out_data_ref <= 8'h3c;
      12'd1368 : out_data_ref <= 8'h56;
      12'd1369 : out_data_ref <= 8'h23;
      12'd1370 : out_data_ref <= 8'h67;
      12'd1371 : out_data_ref <= 8'h74;
      12'd1372 : out_data_ref <= 8'h3d;
      12'd1373 : out_data_ref <= 8'hcd;
      12'd1374 : out_data_ref <= 8'h6e;
      12'd1375 : out_data_ref <= 8'h40;
      12'd1376 : out_data_ref <= 8'hc0;
      12'd1377 : out_data_ref <= 8'h55;
      12'd1378 : out_data_ref <= 8'hc3;
      12'd1379 : out_data_ref <= 8'h24;
      12'd1380 : out_data_ref <= 8'hc2;
      12'd1381 : out_data_ref <= 8'h72;
      12'd1382 : out_data_ref <= 8'h5a;
      12'd1383 : out_data_ref <= 8'h0d;
      12'd1384 : out_data_ref <= 8'hba;
      12'd1385 : out_data_ref <= 8'haa;
      12'd1386 : out_data_ref <= 8'h75;
      12'd1387 : out_data_ref <= 8'h76;
      12'd1388 : out_data_ref <= 8'h28;
      12'd1389 : out_data_ref <= 8'ha1;
      12'd1390 : out_data_ref <= 8'h20;
      12'd1391 : out_data_ref <= 8'h2b;
      12'd1392 : out_data_ref <= 8'h0b;
      12'd1393 : out_data_ref <= 8'h1c;
      12'd1394 : out_data_ref <= 8'h3c;
      12'd1395 : out_data_ref <= 8'hb7;
      12'd1396 : out_data_ref <= 8'hdf;
      12'd1397 : out_data_ref <= 8'hba;
      12'd1398 : out_data_ref <= 8'h0b;
      12'd1399 : out_data_ref <= 8'h09;
      12'd1400 : out_data_ref <= 8'hcf;
      12'd1401 : out_data_ref <= 8'h53;
      12'd1402 : out_data_ref <= 8'h2f;
      12'd1403 : out_data_ref <= 8'h91;
      12'd1404 : out_data_ref <= 8'h94;
      12'd1405 : out_data_ref <= 8'he5;
      12'd1406 : out_data_ref <= 8'h98;
      12'd1407 : out_data_ref <= 8'h72;
      12'd1408 : out_data_ref <= 8'h40;
      12'd1409 : out_data_ref <= 8'h26;
      12'd1410 : out_data_ref <= 8'h0a;
      12'd1411 : out_data_ref <= 8'h7a;
      12'd1412 : out_data_ref <= 8'h28;
      12'd1413 : out_data_ref <= 8'hde;
      12'd1414 : out_data_ref <= 8'hb9;
      12'd1415 : out_data_ref <= 8'h9d;
      12'd1416 : out_data_ref <= 8'hd3;
      12'd1417 : out_data_ref <= 8'h40;
      12'd1418 : out_data_ref <= 8'h9f;
      12'd1419 : out_data_ref <= 8'h81;
      12'd1420 : out_data_ref <= 8'h7d;
      12'd1421 : out_data_ref <= 8'h5c;
      12'd1422 : out_data_ref <= 8'h06;
      12'd1423 : out_data_ref <= 8'h66;
      12'd1424 : out_data_ref <= 8'he2;
      12'd1425 : out_data_ref <= 8'h48;
      12'd1426 : out_data_ref <= 8'h80;
      12'd1427 : out_data_ref <= 8'h64;
      12'd1428 : out_data_ref <= 8'h2f;
      12'd1429 : out_data_ref <= 8'h0a;
      12'd1430 : out_data_ref <= 8'hbb;
      12'd1431 : out_data_ref <= 8'h92;
      12'd1432 : out_data_ref <= 8'ha9;
      12'd1433 : out_data_ref <= 8'h35;
      12'd1434 : out_data_ref <= 8'h90;
      12'd1435 : out_data_ref <= 8'h02;
      12'd1436 : out_data_ref <= 8'h33;
      12'd1437 : out_data_ref <= 8'h9b;
      12'd1438 : out_data_ref <= 8'hce;
      12'd1439 : out_data_ref <= 8'haa;
      12'd1440 : out_data_ref <= 8'haa;
      12'd1441 : out_data_ref <= 8'h2b;
      12'd1442 : out_data_ref <= 8'haf;
      12'd1443 : out_data_ref <= 8'h2d;
      12'd1444 : out_data_ref <= 8'h27;
      12'd1445 : out_data_ref <= 8'h1f;
      12'd1446 : out_data_ref <= 8'hab;
      12'd1447 : out_data_ref <= 8'h7e;
      12'd1448 : out_data_ref <= 8'h5f;
      12'd1449 : out_data_ref <= 8'h16;
      12'd1450 : out_data_ref <= 8'hae;
      12'd1451 : out_data_ref <= 8'ha3;
      12'd1452 : out_data_ref <= 8'h16;
      12'd1453 : out_data_ref <= 8'hf6;
      12'd1454 : out_data_ref <= 8'ha7;
      12'd1455 : out_data_ref <= 8'hde;
      12'd1456 : out_data_ref <= 8'h17;
      12'd1457 : out_data_ref <= 8'h01;
      12'd1458 : out_data_ref <= 8'h7a;
      12'd1459 : out_data_ref <= 8'h0a;
      12'd1460 : out_data_ref <= 8'h9c;
      12'd1461 : out_data_ref <= 8'h7c;
      12'd1462 : out_data_ref <= 8'h70;
      12'd1463 : out_data_ref <= 8'h28;
      12'd1464 : out_data_ref <= 8'hef;
      12'd1465 : out_data_ref <= 8'h59;
      12'd1466 : out_data_ref <= 8'hd6;
      12'd1467 : out_data_ref <= 8'h0b;
      12'd1468 : out_data_ref <= 8'h52;
      12'd1469 : out_data_ref <= 8'he7;
      12'd1470 : out_data_ref <= 8'h75;
      12'd1471 : out_data_ref <= 8'hb6;
      12'd1472 : out_data_ref <= 8'hcd;
      12'd1473 : out_data_ref <= 8'h24;
      12'd1474 : out_data_ref <= 8'heb;
      12'd1475 : out_data_ref <= 8'h0b;
      12'd1476 : out_data_ref <= 8'h20;
      12'd1477 : out_data_ref <= 8'h13;
      12'd1478 : out_data_ref <= 8'h0e;
      12'd1479 : out_data_ref <= 8'hb3;
      12'd1480 : out_data_ref <= 8'hb6;
      12'd1481 : out_data_ref <= 8'h48;
      12'd1482 : out_data_ref <= 8'hea;
      12'd1483 : out_data_ref <= 8'h3f;
      12'd1484 : out_data_ref <= 8'heb;
      12'd1485 : out_data_ref <= 8'hfe;
      12'd1486 : out_data_ref <= 8'h19;
      12'd1487 : out_data_ref <= 8'hf9;
      12'd1488 : out_data_ref <= 8'h16;
      12'd1489 : out_data_ref <= 8'h41;
      12'd1490 : out_data_ref <= 8'h81;
      12'd1491 : out_data_ref <= 8'h5a;
      12'd1492 : out_data_ref <= 8'hfe;
      12'd1493 : out_data_ref <= 8'h10;
      12'd1494 : out_data_ref <= 8'h1b;
      12'd1495 : out_data_ref <= 8'hc0;
      12'd1496 : out_data_ref <= 8'hf2;
      12'd1497 : out_data_ref <= 8'hf7;
      12'd1498 : out_data_ref <= 8'hae;
      12'd1499 : out_data_ref <= 8'haf;
      12'd1500 : out_data_ref <= 8'h57;
      12'd1501 : out_data_ref <= 8'h7d;
      12'd1502 : out_data_ref <= 8'h98;
      12'd1503 : out_data_ref <= 8'h2b;
      12'd1504 : out_data_ref <= 8'h2f;
      12'd1505 : out_data_ref <= 8'he0;
      12'd1506 : out_data_ref <= 8'h16;
      12'd1507 : out_data_ref <= 8'h10;
      12'd1508 : out_data_ref <= 8'h4f;
      12'd1509 : out_data_ref <= 8'h9e;
      12'd1510 : out_data_ref <= 8'h55;
      12'd1511 : out_data_ref <= 8'h60;
      12'd1512 : out_data_ref <= 8'h92;
      12'd1513 : out_data_ref <= 8'hfa;
      12'd1514 : out_data_ref <= 8'h3d;
      12'd1515 : out_data_ref <= 8'h64;
      12'd1516 : out_data_ref <= 8'h39;
      12'd1517 : out_data_ref <= 8'h28;
      12'd1518 : out_data_ref <= 8'he4;
      12'd1519 : out_data_ref <= 8'hf4;
      12'd1520 : out_data_ref <= 8'heb;
      12'd1521 : out_data_ref <= 8'hc7;
      12'd1522 : out_data_ref <= 8'h58;
      12'd1523 : out_data_ref <= 8'h95;
      12'd1524 : out_data_ref <= 8'heb;
      12'd1525 : out_data_ref <= 8'h33;
      12'd1526 : out_data_ref <= 8'h1e;
      12'd1527 : out_data_ref <= 8'h49;
      12'd1528 : out_data_ref <= 8'h41;
      12'd1529 : out_data_ref <= 8'h67;
      12'd1530 : out_data_ref <= 8'ha3;
      12'd1531 : out_data_ref <= 8'h3b;
      12'd1532 : out_data_ref <= 8'h54;
      12'd1533 : out_data_ref <= 8'h16;
      12'd1534 : out_data_ref <= 8'hc4;
      12'd1535 : out_data_ref <= 8'h12;
      12'd1536 : out_data_ref <= 8'ha7;
      12'd1537 : out_data_ref <= 8'hb5;
      12'd1538 : out_data_ref <= 8'h30;
      12'd1539 : out_data_ref <= 8'h29;
      12'd1540 : out_data_ref <= 8'h88;
      12'd1541 : out_data_ref <= 8'ha5;
      12'd1542 : out_data_ref <= 8'hf9;
      12'd1543 : out_data_ref <= 8'h41;
      12'd1544 : out_data_ref <= 8'h84;
      12'd1545 : out_data_ref <= 8'hf9;
      12'd1546 : out_data_ref <= 8'h12;
      12'd1547 : out_data_ref <= 8'h12;
      12'd1548 : out_data_ref <= 8'h37;
      12'd1549 : out_data_ref <= 8'h7f;
      12'd1550 : out_data_ref <= 8'hb9;
      12'd1551 : out_data_ref <= 8'h2d;
      12'd1552 : out_data_ref <= 8'h92;
      12'd1553 : out_data_ref <= 8'h0b;
      12'd1554 : out_data_ref <= 8'h7f;
      12'd1555 : out_data_ref <= 8'ha7;
      12'd1556 : out_data_ref <= 8'h23;
      12'd1557 : out_data_ref <= 8'h19;
      12'd1558 : out_data_ref <= 8'ha5;
      12'd1559 : out_data_ref <= 8'h69;
      12'd1560 : out_data_ref <= 8'h7f;
      12'd1561 : out_data_ref <= 8'h28;
      12'd1562 : out_data_ref <= 8'hde;
      12'd1563 : out_data_ref <= 8'h00;
      12'd1564 : out_data_ref <= 8'hdc;
      12'd1565 : out_data_ref <= 8'ha5;
      12'd1566 : out_data_ref <= 8'h1d;
      12'd1567 : out_data_ref <= 8'he4;
      12'd1568 : out_data_ref <= 8'h1d;
      12'd1569 : out_data_ref <= 8'h99;
      12'd1570 : out_data_ref <= 8'h12;
      12'd1571 : out_data_ref <= 8'h17;
      12'd1572 : out_data_ref <= 8'hde;
      12'd1573 : out_data_ref <= 8'ha1;
      12'd1574 : out_data_ref <= 8'h45;
      12'd1575 : out_data_ref <= 8'hc0;
      12'd1576 : out_data_ref <= 8'hf2;
      12'd1577 : out_data_ref <= 8'h2a;
      12'd1578 : out_data_ref <= 8'h35;
      12'd1579 : out_data_ref <= 8'h4b;
      12'd1580 : out_data_ref <= 8'hc5;
      12'd1581 : out_data_ref <= 8'hcd;
      12'd1582 : out_data_ref <= 8'hb3;
      12'd1583 : out_data_ref <= 8'h07;
      12'd1584 : out_data_ref <= 8'h95;
      12'd1585 : out_data_ref <= 8'hb3;
      12'd1586 : out_data_ref <= 8'hb9;
      12'd1587 : out_data_ref <= 8'hf8;
      12'd1588 : out_data_ref <= 8'ha5;
      12'd1589 : out_data_ref <= 8'hff;
      12'd1590 : out_data_ref <= 8'h4e;
      12'd1591 : out_data_ref <= 8'h95;
      12'd1592 : out_data_ref <= 8'h91;
      12'd1593 : out_data_ref <= 8'h27;
      12'd1594 : out_data_ref <= 8'h44;
      12'd1595 : out_data_ref <= 8'h64;
      12'd1596 : out_data_ref <= 8'hf7;
      12'd1597 : out_data_ref <= 8'h52;
      12'd1598 : out_data_ref <= 8'h3b;
      12'd1599 : out_data_ref <= 8'he5;
      12'd1600 : out_data_ref <= 8'h6d;
      12'd1601 : out_data_ref <= 8'hee;
      12'd1602 : out_data_ref <= 8'h4c;
      12'd1603 : out_data_ref <= 8'h63;
      12'd1604 : out_data_ref <= 8'h73;
      12'd1605 : out_data_ref <= 8'h11;
      12'd1606 : out_data_ref <= 8'ha5;
      12'd1607 : out_data_ref <= 8'h81;
      12'd1608 : out_data_ref <= 8'h4c;
      12'd1609 : out_data_ref <= 8'hbb;
      12'd1610 : out_data_ref <= 8'h14;
      12'd1611 : out_data_ref <= 8'hcf;
      12'd1612 : out_data_ref <= 8'h1d;
      12'd1613 : out_data_ref <= 8'h70;
      12'd1614 : out_data_ref <= 8'h2b;
      12'd1615 : out_data_ref <= 8'h65;
      12'd1616 : out_data_ref <= 8'h34;
      12'd1617 : out_data_ref <= 8'h3b;
      12'd1618 : out_data_ref <= 8'h30;
      12'd1619 : out_data_ref <= 8'h1f;
      12'd1620 : out_data_ref <= 8'hce;
      12'd1621 : out_data_ref <= 8'h79;
      12'd1622 : out_data_ref <= 8'hb4;
      12'd1623 : out_data_ref <= 8'h95;
      12'd1624 : out_data_ref <= 8'hc9;
      12'd1625 : out_data_ref <= 8'h7d;
      12'd1626 : out_data_ref <= 8'he8;
      12'd1627 : out_data_ref <= 8'hb6;
      12'd1628 : out_data_ref <= 8'h6f;
      12'd1629 : out_data_ref <= 8'hf9;
      12'd1630 : out_data_ref <= 8'h01;
      12'd1631 : out_data_ref <= 8'h32;
      12'd1632 : out_data_ref <= 8'h36;
      12'd1633 : out_data_ref <= 8'h14;
      12'd1634 : out_data_ref <= 8'h4d;
      12'd1635 : out_data_ref <= 8'hd0;
      12'd1636 : out_data_ref <= 8'h72;
      12'd1637 : out_data_ref <= 8'h0b;
      12'd1638 : out_data_ref <= 8'h1c;
      12'd1639 : out_data_ref <= 8'h83;
      12'd1640 : out_data_ref <= 8'h5b;
      12'd1641 : out_data_ref <= 8'h54;
      12'd1642 : out_data_ref <= 8'h9f;
      12'd1643 : out_data_ref <= 8'h9f;
      12'd1644 : out_data_ref <= 8'h62;
      12'd1645 : out_data_ref <= 8'hed;
      12'd1646 : out_data_ref <= 8'h9f;
      12'd1647 : out_data_ref <= 8'he4;
      12'd1648 : out_data_ref <= 8'h1a;
      12'd1649 : out_data_ref <= 8'h7a;
      12'd1650 : out_data_ref <= 8'hee;
      12'd1651 : out_data_ref <= 8'h49;
      12'd1652 : out_data_ref <= 8'h1d;
      12'd1653 : out_data_ref <= 8'hcc;
      12'd1654 : out_data_ref <= 8'hfb;
      12'd1655 : out_data_ref <= 8'hb9;
      12'd1656 : out_data_ref <= 8'he6;
      12'd1657 : out_data_ref <= 8'h89;
      12'd1658 : out_data_ref <= 8'hde;
      12'd1659 : out_data_ref <= 8'he7;
      12'd1660 : out_data_ref <= 8'h19;
      12'd1661 : out_data_ref <= 8'h5b;
      12'd1662 : out_data_ref <= 8'hed;
      12'd1663 : out_data_ref <= 8'hef;
      12'd1664 : out_data_ref <= 8'he1;
      12'd1665 : out_data_ref <= 8'ha6;
      12'd1666 : out_data_ref <= 8'h2b;
      12'd1667 : out_data_ref <= 8'h98;
      12'd1668 : out_data_ref <= 8'h19;
      12'd1669 : out_data_ref <= 8'h2b;
      12'd1670 : out_data_ref <= 8'hb1;
      12'd1671 : out_data_ref <= 8'h3c;
      12'd1672 : out_data_ref <= 8'hba;
      12'd1673 : out_data_ref <= 8'haa;
      12'd1674 : out_data_ref <= 8'h13;
      12'd1675 : out_data_ref <= 8'h7a;
      12'd1676 : out_data_ref <= 8'h87;
      12'd1677 : out_data_ref <= 8'h7e;
      12'd1678 : out_data_ref <= 8'hf7;
      12'd1679 : out_data_ref <= 8'hb1;
      12'd1680 : out_data_ref <= 8'h89;
      12'd1681 : out_data_ref <= 8'h5f;
      12'd1682 : out_data_ref <= 8'he3;
      12'd1683 : out_data_ref <= 8'h1e;
      12'd1684 : out_data_ref <= 8'h99;
      12'd1685 : out_data_ref <= 8'hb8;
      12'd1686 : out_data_ref <= 8'h72;
      12'd1687 : out_data_ref <= 8'h61;
      12'd1688 : out_data_ref <= 8'h47;
      12'd1689 : out_data_ref <= 8'h98;
      12'd1690 : out_data_ref <= 8'h11;
      12'd1691 : out_data_ref <= 8'hd5;
      12'd1692 : out_data_ref <= 8'ha0;
      12'd1693 : out_data_ref <= 8'h36;
      12'd1694 : out_data_ref <= 8'h02;
      12'd1695 : out_data_ref <= 8'h91;
      12'd1696 : out_data_ref <= 8'h26;
      12'd1697 : out_data_ref <= 8'h2f;
      12'd1698 : out_data_ref <= 8'h4f;
      12'd1699 : out_data_ref <= 8'h1d;
      12'd1700 : out_data_ref <= 8'h93;
      12'd1701 : out_data_ref <= 8'h1b;
      12'd1702 : out_data_ref <= 8'hf7;
      12'd1703 : out_data_ref <= 8'h38;
      12'd1704 : out_data_ref <= 8'h84;
      12'd1705 : out_data_ref <= 8'h65;
      12'd1706 : out_data_ref <= 8'hfd;
      12'd1707 : out_data_ref <= 8'hcf;
      12'd1708 : out_data_ref <= 8'h6b;
      12'd1709 : out_data_ref <= 8'hf3;
      12'd1710 : out_data_ref <= 8'h7f;
      12'd1711 : out_data_ref <= 8'h27;
      12'd1712 : out_data_ref <= 8'h1c;
      12'd1713 : out_data_ref <= 8'h15;
      12'd1714 : out_data_ref <= 8'hba;
      12'd1715 : out_data_ref <= 8'h6c;
      12'd1716 : out_data_ref <= 8'hfa;
      12'd1717 : out_data_ref <= 8'h4f;
      12'd1718 : out_data_ref <= 8'h91;
      12'd1719 : out_data_ref <= 8'hda;
      12'd1720 : out_data_ref <= 8'ha5;
      12'd1721 : out_data_ref <= 8'h7d;
      12'd1722 : out_data_ref <= 8'h7b;
      12'd1723 : out_data_ref <= 8'h1e;
      12'd1724 : out_data_ref <= 8'haa;
      12'd1725 : out_data_ref <= 8'h58;
      12'd1726 : out_data_ref <= 8'h21;
      12'd1727 : out_data_ref <= 8'h1e;
      12'd1728 : out_data_ref <= 8'hbe;
      12'd1729 : out_data_ref <= 8'h92;
      12'd1730 : out_data_ref <= 8'h59;
      12'd1731 : out_data_ref <= 8'h3e;
      12'd1732 : out_data_ref <= 8'haa;
      12'd1733 : out_data_ref <= 8'hed;
      12'd1734 : out_data_ref <= 8'h81;
      12'd1735 : out_data_ref <= 8'h34;
      12'd1736 : out_data_ref <= 8'h82;
      12'd1737 : out_data_ref <= 8'h7c;
      12'd1738 : out_data_ref <= 8'h45;
      12'd1739 : out_data_ref <= 8'ha0;
      12'd1740 : out_data_ref <= 8'hed;
      12'd1741 : out_data_ref <= 8'h25;
      12'd1742 : out_data_ref <= 8'h3d;
      12'd1743 : out_data_ref <= 8'h9e;
      12'd1744 : out_data_ref <= 8'h0f;
      12'd1745 : out_data_ref <= 8'h10;
      12'd1746 : out_data_ref <= 8'hdf;
      12'd1747 : out_data_ref <= 8'h96;
      12'd1748 : out_data_ref <= 8'h27;
      12'd1749 : out_data_ref <= 8'h28;
      12'd1750 : out_data_ref <= 8'h62;
      12'd1751 : out_data_ref <= 8'h1e;
      12'd1752 : out_data_ref <= 8'ha6;
      12'd1753 : out_data_ref <= 8'h54;
      12'd1754 : out_data_ref <= 8'hd7;
      12'd1755 : out_data_ref <= 8'hbc;
      12'd1756 : out_data_ref <= 8'had;
      12'd1757 : out_data_ref <= 8'h4e;
      12'd1758 : out_data_ref <= 8'h26;
      12'd1759 : out_data_ref <= 8'hcd;
      12'd1760 : out_data_ref <= 8'hbb;
      12'd1761 : out_data_ref <= 8'hcc;
      12'd1762 : out_data_ref <= 8'hb8;
      12'd1763 : out_data_ref <= 8'h1a;
      12'd1764 : out_data_ref <= 8'he5;
      12'd1765 : out_data_ref <= 8'h48;
      12'd1766 : out_data_ref <= 8'h6a;
      12'd1767 : out_data_ref <= 8'h26;
      12'd1768 : out_data_ref <= 8'h01;
      12'd1769 : out_data_ref <= 8'hca;
      12'd1770 : out_data_ref <= 8'h2f;
      12'd1771 : out_data_ref <= 8'hc2;
      12'd1772 : out_data_ref <= 8'h41;
      12'd1773 : out_data_ref <= 8'h80;
      12'd1774 : out_data_ref <= 8'h1b;
      12'd1775 : out_data_ref <= 8'he7;
      12'd1776 : out_data_ref <= 8'h87;
      12'd1777 : out_data_ref <= 8'he7;
      12'd1778 : out_data_ref <= 8'h51;
      12'd1779 : out_data_ref <= 8'h25;
      12'd1780 : out_data_ref <= 8'ha1;
      12'd1781 : out_data_ref <= 8'h63;
      12'd1782 : out_data_ref <= 8'hc3;
      12'd1783 : out_data_ref <= 8'h2b;
      12'd1784 : out_data_ref <= 8'hf1;
      12'd1785 : out_data_ref <= 8'hb2;
      12'd1786 : out_data_ref <= 8'h91;
      12'd1787 : out_data_ref <= 8'ha2;
      12'd1788 : out_data_ref <= 8'hb3;
      12'd1789 : out_data_ref <= 8'hdb;
      12'd1790 : out_data_ref <= 8'he3;
      12'd1791 : out_data_ref <= 8'hb2;
      12'd1792 : out_data_ref <= 8'ha6;
      12'd1793 : out_data_ref <= 8'h70;
      12'd1794 : out_data_ref <= 8'hf8;
      12'd1795 : out_data_ref <= 8'h8a;
      12'd1796 : out_data_ref <= 8'h55;
      12'd1797 : out_data_ref <= 8'hae;
      12'd1798 : out_data_ref <= 8'h57;
      12'd1799 : out_data_ref <= 8'h73;
      12'd1800 : out_data_ref <= 8'h8f;
      12'd1801 : out_data_ref <= 8'h4a;
      12'd1802 : out_data_ref <= 8'h80;
      12'd1803 : out_data_ref <= 8'h41;
      12'd1804 : out_data_ref <= 8'he4;
      12'd1805 : out_data_ref <= 8'h6f;
      12'd1806 : out_data_ref <= 8'h62;
      12'd1807 : out_data_ref <= 8'h0e;
      12'd1808 : out_data_ref <= 8'h07;
      12'd1809 : out_data_ref <= 8'h74;
      12'd1810 : out_data_ref <= 8'h96;
      12'd1811 : out_data_ref <= 8'hd3;
      12'd1812 : out_data_ref <= 8'hf1;
      12'd1813 : out_data_ref <= 8'hae;
      12'd1814 : out_data_ref <= 8'h05;
      12'd1815 : out_data_ref <= 8'h05;
      12'd1816 : out_data_ref <= 8'h77;
      12'd1817 : out_data_ref <= 8'h46;
      12'd1818 : out_data_ref <= 8'hac;
      12'd1819 : out_data_ref <= 8'hf6;
      12'd1820 : out_data_ref <= 8'h5a;
      12'd1821 : out_data_ref <= 8'h63;
      12'd1822 : out_data_ref <= 8'h9c;
      12'd1823 : out_data_ref <= 8'hf3;
      12'd1824 : out_data_ref <= 8'h6c;
      12'd1825 : out_data_ref <= 8'h55;
      12'd1826 : out_data_ref <= 8'hab;
      12'd1827 : out_data_ref <= 8'h4d;
      12'd1828 : out_data_ref <= 8'hce;
      12'd1829 : out_data_ref <= 8'h9a;
      12'd1830 : out_data_ref <= 8'h79;
      12'd1831 : out_data_ref <= 8'h1c;
      12'd1832 : out_data_ref <= 8'h30;
      12'd1833 : out_data_ref <= 8'hbf;
      12'd1834 : out_data_ref <= 8'h8e;
      12'd1835 : out_data_ref <= 8'hbc;
      12'd1836 : out_data_ref <= 8'h1d;
      12'd1837 : out_data_ref <= 8'h0a;
      12'd1838 : out_data_ref <= 8'ha4;
      12'd1839 : out_data_ref <= 8'h8a;
      12'd1840 : out_data_ref <= 8'h2e;
      12'd1841 : out_data_ref <= 8'h2b;
      12'd1842 : out_data_ref <= 8'h71;
      12'd1843 : out_data_ref <= 8'hbd;
      12'd1844 : out_data_ref <= 8'h29;
      12'd1845 : out_data_ref <= 8'h14;
      12'd1846 : out_data_ref <= 8'hb2;
      12'd1847 : out_data_ref <= 8'h0b;
      12'd1848 : out_data_ref <= 8'hfe;
      12'd1849 : out_data_ref <= 8'ha5;
      12'd1850 : out_data_ref <= 8'h67;
      12'd1851 : out_data_ref <= 8'h39;
      12'd1852 : out_data_ref <= 8'h05;
      12'd1853 : out_data_ref <= 8'h48;
      12'd1854 : out_data_ref <= 8'h2d;
      12'd1855 : out_data_ref <= 8'h9b;
      12'd1856 : out_data_ref <= 8'hd5;
      12'd1857 : out_data_ref <= 8'he7;
      12'd1858 : out_data_ref <= 8'hd6;
      12'd1859 : out_data_ref <= 8'h12;
      12'd1860 : out_data_ref <= 8'h05;
      12'd1861 : out_data_ref <= 8'hfa;
      12'd1862 : out_data_ref <= 8'h34;
      12'd1863 : out_data_ref <= 8'h4f;
      12'd1864 : out_data_ref <= 8'hdd;
      12'd1865 : out_data_ref <= 8'h31;
      12'd1866 : out_data_ref <= 8'h63;
      12'd1867 : out_data_ref <= 8'had;
      12'd1868 : out_data_ref <= 8'h59;
      12'd1869 : out_data_ref <= 8'h2c;
      12'd1870 : out_data_ref <= 8'hca;
      12'd1871 : out_data_ref <= 8'h04;
      12'd1872 : out_data_ref <= 8'ha9;
      12'd1873 : out_data_ref <= 8'h40;
      12'd1874 : out_data_ref <= 8'h03;
      12'd1875 : out_data_ref <= 8'h02;
      12'd1876 : out_data_ref <= 8'h99;
      12'd1877 : out_data_ref <= 8'hc9;
      12'd1878 : out_data_ref <= 8'he7;
      12'd1879 : out_data_ref <= 8'h96;
      12'd1880 : out_data_ref <= 8'h5e;
      12'd1881 : out_data_ref <= 8'hf7;
      12'd1882 : out_data_ref <= 8'hc6;
      12'd1883 : out_data_ref <= 8'h71;
      12'd1884 : out_data_ref <= 8'h0f;
      12'd1885 : out_data_ref <= 8'h90;
      12'd1886 : out_data_ref <= 8'he5;
      12'd1887 : out_data_ref <= 8'h43;
      12'd1888 : out_data_ref <= 8'h91;
      12'd1889 : out_data_ref <= 8'h50;
      12'd1890 : out_data_ref <= 8'h4f;
      12'd1891 : out_data_ref <= 8'ha7;
      12'd1892 : out_data_ref <= 8'ha3;
      12'd1893 : out_data_ref <= 8'hf9;
      12'd1894 : out_data_ref <= 8'h6f;
      12'd1895 : out_data_ref <= 8'h48;
      12'd1896 : out_data_ref <= 8'h18;
      12'd1897 : out_data_ref <= 8'h13;
      12'd1898 : out_data_ref <= 8'ha8;
      12'd1899 : out_data_ref <= 8'h6a;
      12'd1900 : out_data_ref <= 8'h63;
      12'd1901 : out_data_ref <= 8'h4c;
      12'd1902 : out_data_ref <= 8'h12;
      12'd1903 : out_data_ref <= 8'h51;
      12'd1904 : out_data_ref <= 8'h83;
      12'd1905 : out_data_ref <= 8'hfb;
      12'd1906 : out_data_ref <= 8'h82;
      12'd1907 : out_data_ref <= 8'hbd;
      12'd1908 : out_data_ref <= 8'h1a;
      12'd1909 : out_data_ref <= 8'h75;
      12'd1910 : out_data_ref <= 8'h3c;
      12'd1911 : out_data_ref <= 8'h88;
      12'd1912 : out_data_ref <= 8'h1f;
      12'd1913 : out_data_ref <= 8'h9b;
      12'd1914 : out_data_ref <= 8'h6b;
      12'd1915 : out_data_ref <= 8'h92;
      12'd1916 : out_data_ref <= 8'h1b;
      12'd1917 : out_data_ref <= 8'hb2;
      12'd1918 : out_data_ref <= 8'h32;
      12'd1919 : out_data_ref <= 8'h36;
      12'd1920 : out_data_ref <= 8'hbd;
      12'd1921 : out_data_ref <= 8'hab;
      12'd1922 : out_data_ref <= 8'h0a;
      12'd1923 : out_data_ref <= 8'h6a;
      12'd1924 : out_data_ref <= 8'h2c;
      12'd1925 : out_data_ref <= 8'h16;
      12'd1926 : out_data_ref <= 8'hc5;
      12'd1927 : out_data_ref <= 8'h42;
      12'd1928 : out_data_ref <= 8'h1e;
      12'd1929 : out_data_ref <= 8'h72;
      12'd1930 : out_data_ref <= 8'h23;
      12'd1931 : out_data_ref <= 8'h99;
      12'd1932 : out_data_ref <= 8'h30;
      12'd1933 : out_data_ref <= 8'hc5;
      12'd1934 : out_data_ref <= 8'he4;
      12'd1935 : out_data_ref <= 8'h57;
      12'd1936 : out_data_ref <= 8'hd2;
      12'd1937 : out_data_ref <= 8'hcf;
      12'd1938 : out_data_ref <= 8'h72;
      12'd1939 : out_data_ref <= 8'hfd;
      12'd1940 : out_data_ref <= 8'hed;
      12'd1941 : out_data_ref <= 8'h66;
      12'd1942 : out_data_ref <= 8'h3d;
      12'd1943 : out_data_ref <= 8'hff;
      12'd1944 : out_data_ref <= 8'h80;
      12'd1945 : out_data_ref <= 8'hc8;
      12'd1946 : out_data_ref <= 8'h34;
      12'd1947 : out_data_ref <= 8'h31;
      12'd1948 : out_data_ref <= 8'h91;
      12'd1949 : out_data_ref <= 8'hd5;
      12'd1950 : out_data_ref <= 8'h69;
      12'd1951 : out_data_ref <= 8'h87;
      12'd1952 : out_data_ref <= 8'h88;
      12'd1953 : out_data_ref <= 8'h6b;
      12'd1954 : out_data_ref <= 8'hc1;
      12'd1955 : out_data_ref <= 8'h2f;
      12'd1956 : out_data_ref <= 8'h0a;
      12'd1957 : out_data_ref <= 8'h8f;
      12'd1958 : out_data_ref <= 8'hb4;
      12'd1959 : out_data_ref <= 8'hb5;
      12'd1960 : out_data_ref <= 8'hc4;
      12'd1961 : out_data_ref <= 8'hdc;
      12'd1962 : out_data_ref <= 8'h4a;
      12'd1963 : out_data_ref <= 8'h81;
      12'd1964 : out_data_ref <= 8'hb6;
      12'd1965 : out_data_ref <= 8'h00;
      12'd1966 : out_data_ref <= 8'h89;
      12'd1967 : out_data_ref <= 8'h29;
      12'd1968 : out_data_ref <= 8'hd9;
      12'd1969 : out_data_ref <= 8'ha5;
      12'd1970 : out_data_ref <= 8'h8f;
      12'd1971 : out_data_ref <= 8'hec;
      12'd1972 : out_data_ref <= 8'h27;
      12'd1973 : out_data_ref <= 8'h45;
      12'd1974 : out_data_ref <= 8'hac;
      12'd1975 : out_data_ref <= 8'had;
      12'd1976 : out_data_ref <= 8'h93;
      12'd1977 : out_data_ref <= 8'he7;
      12'd1978 : out_data_ref <= 8'h79;
      12'd1979 : out_data_ref <= 8'h76;
      12'd1980 : out_data_ref <= 8'h8a;
      12'd1981 : out_data_ref <= 8'hd7;
      12'd1982 : out_data_ref <= 8'h60;
      12'd1983 : out_data_ref <= 8'h3a;
      12'd1984 : out_data_ref <= 8'h72;
      12'd1985 : out_data_ref <= 8'hf8;
      12'd1986 : out_data_ref <= 8'hc9;
      12'd1987 : out_data_ref <= 8'h2c;
      12'd1988 : out_data_ref <= 8'h47;
      12'd1989 : out_data_ref <= 8'hc7;
      12'd1990 : out_data_ref <= 8'h94;
      12'd1991 : out_data_ref <= 8'h6e;
      12'd1992 : out_data_ref <= 8'hf5;
      12'd1993 : out_data_ref <= 8'h0d;
      12'd1994 : out_data_ref <= 8'h44;
      12'd1995 : out_data_ref <= 8'h8f;
      12'd1996 : out_data_ref <= 8'heb;
      12'd1997 : out_data_ref <= 8'he0;
      12'd1998 : out_data_ref <= 8'hc3;
      12'd1999 : out_data_ref <= 8'hb3;
      12'd2000 : out_data_ref <= 8'h8d;
      12'd2001 : out_data_ref <= 8'h03;
      12'd2002 : out_data_ref <= 8'hd8;
      12'd2003 : out_data_ref <= 8'h3b;
      12'd2004 : out_data_ref <= 8'he4;
      12'd2005 : out_data_ref <= 8'h34;
      12'd2006 : out_data_ref <= 8'hde;
      12'd2007 : out_data_ref <= 8'h88;
      12'd2008 : out_data_ref <= 8'h20;
      12'd2009 : out_data_ref <= 8'h53;
      12'd2010 : out_data_ref <= 8'hf4;
      12'd2011 : out_data_ref <= 8'h2d;
      12'd2012 : out_data_ref <= 8'h98;
      12'd2013 : out_data_ref <= 8'he8;
      12'd2014 : out_data_ref <= 8'hb5;
      12'd2015 : out_data_ref <= 8'h02;
      12'd2016 : out_data_ref <= 8'h1d;
      12'd2017 : out_data_ref <= 8'h41;
      12'd2018 : out_data_ref <= 8'h63;
      12'd2019 : out_data_ref <= 8'h35;
      12'd2020 : out_data_ref <= 8'h40;
      12'd2021 : out_data_ref <= 8'h01;
      12'd2022 : out_data_ref <= 8'h82;
      12'd2023 : out_data_ref <= 8'hdb;
      12'd2024 : out_data_ref <= 8'h95;
      12'd2025 : out_data_ref <= 8'h18;
      12'd2026 : out_data_ref <= 8'hb8;
      12'd2027 : out_data_ref <= 8'h3e;
      12'd2028 : out_data_ref <= 8'hab;
      12'd2029 : out_data_ref <= 8'h47;
      12'd2030 : out_data_ref <= 8'hdd;
      12'd2031 : out_data_ref <= 8'h25;
      12'd2032 : out_data_ref <= 8'h2f;
      12'd2033 : out_data_ref <= 8'h7e;
      12'd2034 : out_data_ref <= 8'h15;
      12'd2035 : out_data_ref <= 8'hdf;
      12'd2036 : out_data_ref <= 8'h0c;
      12'd2037 : out_data_ref <= 8'h13;
      12'd2038 : out_data_ref <= 8'h91;
      12'd2039 : out_data_ref <= 8'h08;
      12'd2040 : out_data_ref <= 8'h2c;
      12'd2041 : out_data_ref <= 8'h6b;
      12'd2042 : out_data_ref <= 8'h90;
      12'd2043 : out_data_ref <= 8'ha5;
      12'd2044 : out_data_ref <= 8'hfc;
      12'd2045 : out_data_ref <= 8'h10;
      12'd2046 : out_data_ref <= 8'hb8;
      12'd2047 : out_data_ref <= 8'h87;
      12'd2048 : out_data_ref <= 8'h48;
      12'd2049 : out_data_ref <= 8'hf7;
      12'd2050 : out_data_ref <= 8'h78;
      12'd2051 : out_data_ref <= 8'h8c;
      12'd2052 : out_data_ref <= 8'h46;
      12'd2053 : out_data_ref <= 8'h85;
      12'd2054 : out_data_ref <= 8'he7;
      12'd2055 : out_data_ref <= 8'h25;
      12'd2056 : out_data_ref <= 8'h0b;
      12'd2057 : out_data_ref <= 8'h9d;
      12'd2058 : out_data_ref <= 8'h21;
      12'd2059 : out_data_ref <= 8'hde;
      12'd2060 : out_data_ref <= 8'h75;
      12'd2061 : out_data_ref <= 8'h23;
      12'd2062 : out_data_ref <= 8'hdf;
      12'd2063 : out_data_ref <= 8'hf3;
      12'd2064 : out_data_ref <= 8'h7a;
      12'd2065 : out_data_ref <= 8'hae;
      12'd2066 : out_data_ref <= 8'h0a;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
