module ntt16384_163841 ( clk, rst, start, input_fg, addr, din, dout, valid );

  localparam Q0 = 163841;

  // STATE
  localparam ST_IDLE   = 0;
  localparam ST_NTT    = 1;
  localparam ST_PMUL   = 2;
  localparam ST_RELOAD = 3;
  localparam ST_INTT   = 4;
  localparam ST_CRT    = 5;  // not applied for single prime scheme
  localparam ST_REDUCE = 6;
  localparam ST_FINISH = 7;

  input                      clk;
  input                      rst;
  input                      start;
  input                      input_fg;
  input             [14 : 0] addr;
  input signed      [17 : 0] din;
  output reg signed [17 : 0] dout;
  output reg                 valid;

  // BRAM
  reg            wr_en   [0 : 1];
  reg   [14 : 0] wr_addr [0 : 1];
  reg   [14 : 0] rd_addr [0 : 1];
  reg   [17 : 0] wr_din  [0 : 1];
  wire  [17 : 0] rd_dout [0 : 1];
  wire  [17 : 0] wr_dout [0 : 1];

  // addr_gen
  wire         bank_index_rd [0 : 1];
  wire         bank_index_wr [0 : 1];
  wire [13: 0] data_index_rd [0 : 1];
  wire [13: 0] data_index_wr [0 : 1];
  reg  bank_index_wr_0_shift_1, bank_index_wr_0_shift_2;
  reg  fg_shift_1, fg_shift_2, fg_shift_3;

  // w_addr_gen
  reg  [13 : 0] stage_bit;
  wire [13 : 0] w_addr;

  // bfu
  reg                  ntt_state; 
  reg  signed [17: 0] in_a  ;
  reg  signed [17: 0] in_b  ;
  reg  signed [17: 0] in_w  ;
  wire signed [35: 0] bw    ;
  wire signed [17: 0] out_a ;
  wire signed [17: 0] out_b ;

  // state, stage, counter
  reg  [2 : 0] state, next_state;
  reg  [4 : 0] stage, stage_wr;
  wire [4 : 0] stage_rdM, stage_wrM;
  reg  [15 : 0] ctr;
  reg  [15 : 0] ctr_shift_7, ctr_shift_8, ctr_shift_9, ctr_shift_1, ctr_shift_2;
  reg          ctr_MSB_masked;
  reg          poly_select;
  reg          ctr_msb_shift_1;
  wire         ctr_half_end, ctr_full_end, ctr_shift_7_end, stage_rd_end, stage_rd_2, stage_wr_end, ntt_end, point_proc_end, reduce_end;

  // w_array
  reg         [14: 0] w_addr_in;
  wire signed [17: 0] w_dout ;

  // misc
  reg          bank_index_rd_shift_1, bank_index_rd_shift_2;
  reg [14: 0] wr_ctr [0 : 1];
  reg [17: 0] din_shift_1, din_shift_2, din_shift_3;
  reg [14: 0] w_addr_in_shift_1;

  // BRAM instances
  bram_18_15_P bank_0
  (clk, wr_en[0], wr_addr[0], rd_addr[0], wr_din[0], wr_dout[0], rd_dout[0]);
  bram_18_15_P bank_1
  (clk, wr_en[1], wr_addr[1], rd_addr[1], wr_din[1], wr_dout[1], rd_dout[1]);

  // Read/Write Address Generator
  addr_gen addr_rd_0 (clk, stage_rdM, {ctr_MSB_masked, ctr[13:0]}, bank_index_rd[0], data_index_rd[0]);
  addr_gen addr_rd_1 (clk, stage_rdM, {1'b1, ctr[13:0]}, bank_index_rd[1], data_index_rd[1]);
  addr_gen addr_wr_0 (clk, stage_wrM, {wr_ctr[0]}, bank_index_wr[0], data_index_wr[0]);
  addr_gen addr_wr_1 (clk, stage_wrM, {wr_ctr[1]}, bank_index_wr[1], data_index_wr[1]);

  // Omega Address Generator
  w_addr_gen w_addr_gen_0 (clk, stage_bit, ctr[13:0], w_addr);

  // Butterfly Unit  , each with a corresponding omega array
  bfu_163841 bfu_inst (clk, ntt_state, in_a, in_b, in_w, bw, out_a, out_b);
  w_163841 rom_w_inst (clk, w_addr_in_shift_1, w_dout);

  assign ctr_half_end         = (ctr[13:0] == 16383) ? 1 : 0;
  assign ctr_full_end         = (ctr[14:0] == 32767) ? 1 : 0;
  assign stage_rd_end         = (stage == 15) ? 1 : 0;
  assign stage_rd_2           = (stage == 2) ? 1 : 0;
  assign ntt_end         = (stage_rd_end && ctr[13 : 0] == 10) ? 1 : 0;
  assign crt_end         = (stage_rd_2 && ctr[13 : 0] == 10) ? 1 : 0;
  assign point_proc_end   = (ctr == 32778) ? 1 : 0;
  assign reload_end      = (stage != 0 && ctr[13:0] == 4) ? 1 : 0;
  assign reduce_end      = (ctr == 32772);

  // crt
  // fg_shift
  always @ ( posedge clk ) begin
    fg_shift_1 <= input_fg;
    fg_shift_2 <= fg_shift_1;
    fg_shift_3 <= fg_shift_2;
  end
  // dout
  always @ ( posedge clk ) begin
    if (state == ST_FINISH) begin
      if (bank_index_wr_0_shift_2) begin
        dout <= wr_dout[1][17:0];
      end else begin
        dout <= wr_dout[0][17:0];
      end
    end else begin
      dout <= 'sd0;
    end
  end

  // bank_index_wr_0_shift_1
  always @ ( posedge clk ) begin
    bank_index_wr_0_shift_1 <= bank_index_wr[0];
    bank_index_wr_0_shift_2 <= bank_index_wr_0_shift_1;
  end

  // poly_select
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        poly_select <= ~poly_select;
      end else begin
        poly_select <= poly_select;
      end    
    end else if (state == ST_RELOAD) begin
      poly_select <= 1;
    end else begin
      poly_select <= 0;
    end
  end

  // w_addr_in_shift_1
  always @ ( posedge clk ) begin
    w_addr_in_shift_1 <= w_addr_in;
  end

  // din_shift
  always @ ( posedge clk ) begin
    din_shift_1 <= din;
    din_shift_2 <= din_shift_1;
    din_shift_3 <= din_shift_2;
  end

  // rd_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_rd[0]) begin
        rd_addr[0][13:0] <= data_index_rd[1];
        rd_addr[1][13:0] <= data_index_rd[0];
      end else begin
        rd_addr[0][13:0] <= data_index_rd[0];
        rd_addr[1][13:0] <= data_index_rd[1];
      end
    end else begin
      rd_addr[0][13:0] <= data_index_rd[0];
      rd_addr[1][13:0] <= data_index_rd[0];
    end

    if (state == ST_NTT)  begin
      rd_addr[0][14] <= poly_select;
      rd_addr[1][14] <= poly_select;
    end else if (state == ST_PMUL) begin
      rd_addr[0][14] <=  bank_index_rd[0];
      rd_addr[1][14] <= ~bank_index_rd[0];
    end else if (state == ST_RELOAD) begin
      rd_addr[0][14] <= 0;
      rd_addr[1][14] <= 0;
    end else begin
      rd_addr[0][14] <= 1;
      rd_addr[1][14] <= 1;
    end
  end

  // wr_en
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 1;
      end
    end else if (state == ST_IDLE) begin
      if (fg_shift_3 ^ bank_index_wr[0]) begin
        wr_en[0] <= 0;
        wr_en[1] <= 1;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 0;
      end
    end else if (state == ST_PMUL) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_REDUCE) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_CRT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else if (state == ST_RELOAD) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else begin
      wr_en[0] <= 0;
      wr_en[1] <= 0;
    end
  end

  // wr_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_addr[0][13:0] <= data_index_wr[1];
        wr_addr[1][13:0] <= data_index_wr[0];
      end else begin
        wr_addr[0][13:0] <= data_index_wr[0];
        wr_addr[1][13:0] <= data_index_wr[1];
      end
    end else begin
      wr_addr[0][13:0] <= data_index_wr[0];
      wr_addr[1][13:0] <= data_index_wr[0];
    end  

    if (state == ST_IDLE) begin
      wr_addr[0][14] <= fg_shift_3;
      wr_addr[1][14] <= fg_shift_3;
    end else if(state == ST_NTT || state == ST_INTT) begin
      wr_addr[0][14] <= poly_select;
      wr_addr[1][14] <= poly_select;
    end else if (state == ST_PMUL || state == ST_REDUCE || state == ST_FINISH) begin
      wr_addr[0][14] <= 0;
      wr_addr[1][14] <= 0;
    end else begin
      wr_addr[0][14] <= 1;
      wr_addr[1][14] <= 1;
    end     
  end

  // wr_din
  always @ ( posedge clk ) begin
    if (state == ST_IDLE) begin
      wr_din[0][17:0] <= { din_shift_3 };
      wr_din[1][17:0] <= { din_shift_3 };
    end else if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_din[0][17:0] <= out_b;
        wr_din[1][17:0] <= out_a;
      end else begin
        wr_din[0][17:0] <= out_a;
        wr_din[1][17:0] <= out_b;
      end
    end else if (state == ST_RELOAD) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end
    end else if (state == ST_REDUCE) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end
    end else begin
      wr_din[0][17:0] <= out_a;
      wr_din[1][17:0] <= out_a;
    end
  end

  // bank_index_rd_shift
  always @ ( posedge clk ) begin
    bank_index_rd_shift_1 <= bank_index_rd[0];
    bank_index_rd_shift_2 <= bank_index_rd_shift_1;
  end

  // ntt_state
  always @ ( posedge clk ) begin
    if (state == ST_INTT) begin
      ntt_state <= 1;
    end else begin
      ntt_state <= 0;
    end
  end

  // in_a, in_b
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else if (state == ST_CRT) begin
      if (bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else begin // ST_PMUL
      in_b <= $signed(rd_dout[1]);
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_a <= $signed(rd_dout[1]);
      end else begin
        in_a <= $signed(rd_dout[0]);
      end
    end else begin // ST_PMUL, ST_CRT
      in_a <= 'sd0;
    end
  end

  // w_addr_in, in_w
  always @ ( posedge clk ) begin
    if (state == ST_NTT) begin
      w_addr_in <= {1'b0, w_addr};
    end else begin
      w_addr_in <= 32768 - w_addr;
    end

    if (state == ST_PMUL) begin
        in_w <= rd_dout[0];
    end else begin
      in_w <= w_dout;
    end
  end

  // wr_ctr
  always @ ( posedge clk ) begin
    if (state == ST_IDLE || state == ST_FINISH) begin
      wr_ctr[0] <= addr[14:0];
    end else if (state == ST_RELOAD || state == ST_REDUCE) begin
      wr_ctr[0] <= {ctr_shift_1[0], ctr_shift_1[1], ctr_shift_1[2], ctr_shift_1[3], ctr_shift_1[4], ctr_shift_1[5], ctr_shift_1[6], ctr_shift_1[7], ctr_shift_1[8], ctr_shift_1[9], ctr_shift_1[10], ctr_shift_1[11], ctr_shift_1[12], ctr_shift_1[13], ctr_shift_1[14]};
    end else if (state == ST_NTT || state == ST_INTT) begin
      wr_ctr[0] <= {1'b0, ctr_shift_7[13:0]};
    end else begin
      wr_ctr[0] <= ctr_shift_7[14:0];
    end

    wr_ctr[1] <= {1'b1, ctr_shift_7[13:0]};
  end

  // ctr_MSB_masked
  always @ (*) begin
    if (state == ST_NTT || state == ST_INTT) begin
      ctr_MSB_masked = 0;
    end else begin
      ctr_MSB_masked = ctr[14];
    end
  end

  // ctr, ctr_shifts
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_PMUL) begin
      if (point_proc_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_CRT) begin
      if (crt_end || ctr_full_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_REDUCE) begin
      if (reduce_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else begin
      ctr <= 0;
    end

    //change ctr_shift_7 <= ctr - 5;
    ctr_shift_7 <= ctr - 7;
    ctr_shift_8 <= ctr_shift_7;
    ctr_shift_9 <= ctr_shift_8;
    ctr_shift_1 <= ctr;
    ctr_shift_2 <= ctr_shift_1;
  end

  // stage, stage_wr
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage <= 0;
      end else if (ctr_half_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else begin
      stage <= 0;
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[13:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[14:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_9[14:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else begin
      stage_wr <= 0;
    end        
  end
  assign stage_rdM = (state == ST_NTT || state == ST_INTT) ? stage : 0;
  assign stage_wrM = (state == ST_NTT || state == ST_INTT) ? stage_wr : 0;

  // stage_bit
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_bit <= 0;
      end else if (ctr_half_end) begin
        stage_bit[0] <= 1'b1;
        stage_bit[13 : 1] <= stage_bit[12 : 0];
      end else begin
        stage_bit <= stage_bit;
      end
    end else begin
      stage_bit <= 'b0;
    end
  end

  // valid
  always @ (*) begin
      if (state == ST_FINISH) begin
          valid = 1;
      end else begin
          valid = 0;
      end
  end

  // state
  always @ ( posedge clk ) begin
    if(rst) begin
            state <= 0;
        end else begin
            state <= next_state;
        end
  end

  always @(*) begin
    case(state)
    ST_IDLE: begin
      if(start)
        next_state = ST_NTT;
      else
        next_state = ST_IDLE;
    end
    ST_NTT: begin
      if(ntt_end && poly_select == 1)
        next_state = ST_PMUL;
      else
        next_state = ST_NTT;
    end
    ST_PMUL: begin
      if (point_proc_end)
        next_state = ST_RELOAD;
      else
        next_state = ST_PMUL;
    end
    ST_RELOAD: begin
      if (reload_end) begin
        next_state = ST_INTT;
      end else begin
        next_state = ST_RELOAD;
      end
    end
    ST_INTT: begin
      if(ntt_end)
        next_state = ST_REDUCE;
      else
        next_state = ST_INTT;
      end
    ST_REDUCE: begin
      if(reduce_end)
        next_state = ST_FINISH;
      else
        next_state = ST_REDUCE;
    end
    ST_FINISH: begin
      if(!start)
        next_state = ST_FINISH;
      else
        next_state = ST_IDLE;
    end
    default: next_state = ST_IDLE;
    endcase
  end

endmodule

module w_addr_gen ( clk, stage_bit, ctr, w_addr );

  input              clk;
  input      [13: 0] stage_bit;
  input      [13: 0] ctr;
  output reg [13: 0] w_addr;

  wire [13: 0] w;

  assign w[ 0] = (stage_bit[ 0]) ? ctr[ 0] : 0;
  assign w[ 1] = (stage_bit[ 1]) ? ctr[ 1] : 0;
  assign w[ 2] = (stage_bit[ 2]) ? ctr[ 2] : 0;
  assign w[ 3] = (stage_bit[ 3]) ? ctr[ 3] : 0;
  assign w[ 4] = (stage_bit[ 4]) ? ctr[ 4] : 0;
  assign w[ 5] = (stage_bit[ 5]) ? ctr[ 5] : 0;
  assign w[ 6] = (stage_bit[ 6]) ? ctr[ 6] : 0;
  assign w[ 7] = (stage_bit[ 7]) ? ctr[ 7] : 0;
  assign w[ 8] = (stage_bit[ 8]) ? ctr[ 8] : 0;
  assign w[ 9] = (stage_bit[ 9]) ? ctr[ 9] : 0;
  assign w[10] = (stage_bit[10]) ? ctr[10] : 0;
  assign w[11] = (stage_bit[11]) ? ctr[11] : 0;
  assign w[12] = (stage_bit[12]) ? ctr[12] : 0;
  assign w[13] = (stage_bit[13]) ? ctr[13] : 0;

  always @ ( posedge clk ) begin
    w_addr <= {w[0], w[1], w[2], w[3], w[4], w[5], w[6], w[7], w[8], w[9], w[10], w[11], w[12], w[13]};
  end

endmodule

module addr_gen ( clk, stage, ctr, bank_index, data_index );

  input              clk;
  input      [3 : 0] stage;
  input      [14: 0] ctr;
  output reg         bank_index;
  output reg [13: 0] data_index;

  wire       [14: 0] bs_out;

  barrel_shifter bs ( clk, ctr, stage, bs_out );

    always @( posedge clk ) begin
        bank_index <= ^bs_out;
    end

    always @( posedge clk ) begin
        data_index <= bs_out[14:1];
    end

endmodule

module barrel_shifter ( clk, in, shift, out );

  input              clk;
  input      [14: 0] in;
  input      [3 : 0] shift;
  output reg [14: 0] out;

  reg        [14: 0] in_s [0:4];

  always @ (*) begin
    in_s[0] = in;
  end

  always @ (*) begin
    if(shift[0]) begin
      in_s[1] = { in_s[0][0], in_s[0][14:1] };
    end else begin
      in_s[1] = in_s[0];
    end
  end

  always @ (*) begin
    if(shift[1]) begin
      in_s[2] = { in_s[1][1:0], in_s[1][14:2] };
    end else begin
      in_s[2] = in_s[1];
    end
  end

  always @ (*) begin
    if(shift[2]) begin
      in_s[3] = { in_s[2][3:0], in_s[2][14:4] };
    end else begin
      in_s[3] = in_s[2];
    end
  end

  always @ (*) begin
    if(shift[3]) begin
      in_s[4] = { in_s[3][7:0], in_s[3][14:8] };
    end else begin
      in_s[4] = in_s[3];
    end
  end

  always @ ( posedge clk ) begin
    out <= in_s[4];
  end

endmodule

module bfu_163841 ( clk, state, in_a, in_b, w, bw, out_a, out_b );

  input                      clk;
  input                      state;
  input      signed [17 : 0] in_a;
  input      signed [17 : 0] in_b;
  input      signed [17 : 0] w;
  output reg signed [34 : 0] bw;
  output reg signed [17 : 0] out_a;
  output reg signed [17 : 0] out_b;

  wire signed       [17 : 0] mod_bw;
  reg signed        [18 : 0] a, b;
  reg signed        [17 : 0] in_a_s1, in_a_s2, in_a_s3, in_a_s4, in_a_s5;

  reg signed        [34 : 0] bwQ_0, bwQ_1, bwQ_2;
  wire signed       [18 : 0] a_add_q, a_sub_q, b_add_q, b_sub_q;

  modmul163841s mod163841s_inst ( clk, 1'b0, bw, mod_bw );

  assign a_add_q = a + 'sd163841;
  assign a_sub_q = a - 'sd163841;
  assign b_add_q = b + 'sd163841;
  assign b_sub_q = b - 'sd163841;

  always @(posedge clk ) begin
    in_a_s1 <= in_a;
    in_a_s2 <= in_a_s1;
    in_a_s3 <= in_a_s2;
    in_a_s4 <= in_a_s3;
    in_a_s5 <= in_a_s4;
  end

  always @ ( posedge clk ) begin
    bw <= in_b * w;
  end

  always @ ( posedge clk ) begin
    a <= in_a_s4 + mod_bw;
    b <= in_a_s4 - mod_bw;

    if (state == 0) begin
      if (a > 'sd81920) begin
        out_a <= a_sub_q;
      end else if (a < -'sd81920) begin
        out_a <= a_add_q;
      end else begin
        out_a <= a;
      end
    end else begin
      if (a[0] == 0) begin
        out_a <= a[18:1];
      end else if (a[18] == 0) begin // a > 0
        out_a <= a_sub_q[18:1];
      end else begin                 // a < 0
        out_a <= a_add_q[18:1];
      end
    end

    if (state == 0) begin
      if (b > 'sd81920) begin
        out_b <= b_sub_q;
      end else if (b < -'sd81920) begin
        out_b <= b_add_q;
      end else begin
        out_b <= b;
      end
    end else begin
      if (b[0] == 0) begin
        out_b <= b[18:1];
      end else if (b[18] == 0) begin // b > 0
        out_b <= b_sub_q[18:1];
      end else begin                 // b < 0
        out_b <= b_add_q[18:1];
      end
    end
  end

endmodule

module w_163841 ( clk, addr, dout );

  input                       clk;
  input             [14 : 0]  addr;
  output signed     [17 : 0]  dout;

  wire signed       [17 : 0]  dout_p;
  wire signed       [17 : 0]  dout_n;
  reg               [14 : 0]  addr_reg;

  (* rom_style = "block" *) reg signed [17:0] data [0:16383];

  assign dout_p = data[addr_reg[13:0]];
  assign dout_n = -dout_p;
  assign dout   = addr_reg[14] ? dout_n : dout_p;

  always @ ( posedge clk ) begin
    addr_reg <= addr;
  end

  initial begin
    data[    0] =  'sd1;
    data[    1] =  'sd7;
    data[    2] =  'sd49;
    data[    3] =  'sd343;
    data[    4] =  'sd2401;
    data[    5] =  'sd16807;
    data[    6] = -'sd46192;
    data[    7] =  'sd4338;
    data[    8] =  'sd30366;
    data[    9] =  'sd48721;
    data[   10] =  'sd13365;
    data[   11] = -'sd70286;
    data[   12] = -'sd479;
    data[   13] = -'sd3353;
    data[   14] = -'sd23471;
    data[   15] = -'sd456;
    data[   16] = -'sd3192;
    data[   17] = -'sd22344;
    data[   18] =  'sd7433;
    data[   19] =  'sd52031;
    data[   20] =  'sd36535;
    data[   21] = -'sd71937;
    data[   22] = -'sd12036;
    data[   23] =  'sd79589;
    data[   24] =  'sd65600;
    data[   25] = -'sd32323;
    data[   26] = -'sd62420;
    data[   27] =  'sd54583;
    data[   28] =  'sd54399;
    data[   29] =  'sd53111;
    data[   30] =  'sd44095;
    data[   31] = -'sd19017;
    data[   32] =  'sd30722;
    data[   33] =  'sd51213;
    data[   34] =  'sd30809;
    data[   35] =  'sd51822;
    data[   36] =  'sd35072;
    data[   37] =  'sd81663;
    data[   38] =  'sd80118;
    data[   39] =  'sd69303;
    data[   40] = -'sd6402;
    data[   41] = -'sd44814;
    data[   42] =  'sd13984;
    data[   43] = -'sd65953;
    data[   44] =  'sd29852;
    data[   45] =  'sd45123;
    data[   46] = -'sd11821;
    data[   47] =  'sd81094;
    data[   48] =  'sd76135;
    data[   49] =  'sd41422;
    data[   50] = -'sd37728;
    data[   51] =  'sd63586;
    data[   52] = -'sd46421;
    data[   53] =  'sd2735;
    data[   54] =  'sd19145;
    data[   55] = -'sd29826;
    data[   56] = -'sd44941;
    data[   57] =  'sd13095;
    data[   58] = -'sd72176;
    data[   59] = -'sd13709;
    data[   60] =  'sd67878;
    data[   61] = -'sd16377;
    data[   62] =  'sd49202;
    data[   63] =  'sd16732;
    data[   64] = -'sd46717;
    data[   65] =  'sd663;
    data[   66] =  'sd4641;
    data[   67] =  'sd32487;
    data[   68] =  'sd63568;
    data[   69] = -'sd46547;
    data[   70] =  'sd1853;
    data[   71] =  'sd12971;
    data[   72] = -'sd73044;
    data[   73] = -'sd19785;
    data[   74] =  'sd25346;
    data[   75] =  'sd13581;
    data[   76] = -'sd68774;
    data[   77] =  'sd10105;
    data[   78] =  'sd70735;
    data[   79] =  'sd3622;
    data[   80] =  'sd25354;
    data[   81] =  'sd13637;
    data[   82] = -'sd68382;
    data[   83] =  'sd12849;
    data[   84] = -'sd73898;
    data[   85] = -'sd25763;
    data[   86] = -'sd16500;
    data[   87] =  'sd48341;
    data[   88] =  'sd10705;
    data[   89] =  'sd74935;
    data[   90] =  'sd33022;
    data[   91] =  'sd67313;
    data[   92] = -'sd20332;
    data[   93] =  'sd21517;
    data[   94] = -'sd13222;
    data[   95] =  'sd71287;
    data[   96] =  'sd7486;
    data[   97] =  'sd52402;
    data[   98] =  'sd39132;
    data[   99] = -'sd53758;
    data[  100] = -'sd48624;
    data[  101] = -'sd12686;
    data[  102] =  'sd75039;
    data[  103] =  'sd33750;
    data[  104] =  'sd72409;
    data[  105] =  'sd15340;
    data[  106] = -'sd56461;
    data[  107] = -'sd67545;
    data[  108] =  'sd18708;
    data[  109] = -'sd32885;
    data[  110] = -'sd66354;
    data[  111] =  'sd27045;
    data[  112] =  'sd25474;
    data[  113] =  'sd14477;
    data[  114] = -'sd62502;
    data[  115] =  'sd54009;
    data[  116] =  'sd50381;
    data[  117] =  'sd24985;
    data[  118] =  'sd11054;
    data[  119] =  'sd77378;
    data[  120] =  'sd50123;
    data[  121] =  'sd23179;
    data[  122] = -'sd1588;
    data[  123] = -'sd11116;
    data[  124] = -'sd77812;
    data[  125] = -'sd53161;
    data[  126] = -'sd44445;
    data[  127] =  'sd16567;
    data[  128] = -'sd47872;
    data[  129] = -'sd7422;
    data[  130] = -'sd51954;
    data[  131] = -'sd35996;
    data[  132] =  'sd75710;
    data[  133] =  'sd38447;
    data[  134] = -'sd58553;
    data[  135] =  'sd81652;
    data[  136] =  'sd80041;
    data[  137] =  'sd68764;
    data[  138] = -'sd10175;
    data[  139] = -'sd71225;
    data[  140] = -'sd7052;
    data[  141] = -'sd49364;
    data[  142] = -'sd17866;
    data[  143] =  'sd38779;
    data[  144] = -'sd56229;
    data[  145] = -'sd65921;
    data[  146] =  'sd30076;
    data[  147] =  'sd46691;
    data[  148] = -'sd845;
    data[  149] = -'sd5915;
    data[  150] = -'sd41405;
    data[  151] =  'sd37847;
    data[  152] = -'sd62753;
    data[  153] =  'sd52252;
    data[  154] =  'sd38082;
    data[  155] = -'sd61108;
    data[  156] =  'sd63767;
    data[  157] = -'sd45154;
    data[  158] =  'sd11604;
    data[  159] =  'sd81228;
    data[  160] =  'sd77073;
    data[  161] =  'sd47988;
    data[  162] =  'sd8234;
    data[  163] =  'sd57638;
    data[  164] =  'sd75784;
    data[  165] =  'sd38965;
    data[  166] = -'sd54927;
    data[  167] = -'sd56807;
    data[  168] = -'sd69967;
    data[  169] =  'sd1754;
    data[  170] =  'sd12278;
    data[  171] = -'sd77895;
    data[  172] = -'sd53742;
    data[  173] = -'sd48512;
    data[  174] = -'sd11902;
    data[  175] =  'sd80527;
    data[  176] =  'sd72166;
    data[  177] =  'sd13639;
    data[  178] = -'sd68368;
    data[  179] =  'sd12947;
    data[  180] = -'sd73212;
    data[  181] = -'sd20961;
    data[  182] =  'sd17114;
    data[  183] = -'sd44043;
    data[  184] =  'sd19381;
    data[  185] = -'sd28174;
    data[  186] = -'sd33377;
    data[  187] = -'sd69798;
    data[  188] =  'sd2937;
    data[  189] =  'sd20559;
    data[  190] = -'sd19928;
    data[  191] =  'sd24345;
    data[  192] =  'sd6574;
    data[  193] =  'sd46018;
    data[  194] = -'sd5556;
    data[  195] = -'sd38892;
    data[  196] =  'sd55438;
    data[  197] =  'sd60384;
    data[  198] = -'sd68835;
    data[  199] =  'sd9678;
    data[  200] =  'sd67746;
    data[  201] = -'sd17301;
    data[  202] =  'sd42734;
    data[  203] = -'sd28544;
    data[  204] = -'sd35967;
    data[  205] =  'sd75913;
    data[  206] =  'sd39868;
    data[  207] = -'sd48606;
    data[  208] = -'sd12560;
    data[  209] =  'sd75921;
    data[  210] =  'sd39924;
    data[  211] = -'sd48214;
    data[  212] = -'sd9816;
    data[  213] = -'sd68712;
    data[  214] =  'sd10539;
    data[  215] =  'sd73773;
    data[  216] =  'sd24888;
    data[  217] =  'sd10375;
    data[  218] =  'sd72625;
    data[  219] =  'sd16852;
    data[  220] = -'sd45877;
    data[  221] =  'sd6543;
    data[  222] =  'sd45801;
    data[  223] = -'sd7075;
    data[  224] = -'sd49525;
    data[  225] = -'sd18993;
    data[  226] =  'sd30890;
    data[  227] =  'sd52389;
    data[  228] =  'sd39041;
    data[  229] = -'sd54395;
    data[  230] = -'sd53083;
    data[  231] = -'sd43899;
    data[  232] =  'sd20389;
    data[  233] = -'sd21118;
    data[  234] =  'sd16015;
    data[  235] = -'sd51736;
    data[  236] = -'sd34470;
    data[  237] = -'sd77449;
    data[  238] = -'sd50620;
    data[  239] = -'sd26658;
    data[  240] = -'sd22765;
    data[  241] =  'sd4486;
    data[  242] =  'sd31402;
    data[  243] =  'sd55973;
    data[  244] =  'sd64129;
    data[  245] = -'sd42620;
    data[  246] =  'sd29342;
    data[  247] =  'sd41553;
    data[  248] = -'sd36811;
    data[  249] =  'sd70005;
    data[  250] = -'sd1488;
    data[  251] = -'sd10416;
    data[  252] = -'sd72912;
    data[  253] = -'sd18861;
    data[  254] =  'sd31814;
    data[  255] =  'sd58857;
    data[  256] = -'sd79524;
    data[  257] = -'sd65145;
    data[  258] =  'sd35508;
    data[  259] = -'sd79126;
    data[  260] = -'sd62359;
    data[  261] =  'sd55010;
    data[  262] =  'sd57388;
    data[  263] =  'sd74034;
    data[  264] =  'sd26715;
    data[  265] =  'sd23164;
    data[  266] = -'sd1693;
    data[  267] = -'sd11851;
    data[  268] =  'sd80884;
    data[  269] =  'sd74665;
    data[  270] =  'sd31132;
    data[  271] =  'sd54083;
    data[  272] =  'sd50899;
    data[  273] =  'sd28611;
    data[  274] =  'sd36436;
    data[  275] = -'sd72630;
    data[  276] = -'sd16887;
    data[  277] =  'sd45632;
    data[  278] = -'sd8258;
    data[  279] = -'sd57806;
    data[  280] = -'sd76960;
    data[  281] = -'sd47197;
    data[  282] = -'sd2697;
    data[  283] = -'sd18879;
    data[  284] =  'sd31688;
    data[  285] =  'sd57975;
    data[  286] =  'sd78143;
    data[  287] =  'sd55478;
    data[  288] =  'sd60664;
    data[  289] = -'sd66875;
    data[  290] =  'sd23398;
    data[  291] = -'sd55;
    data[  292] = -'sd385;
    data[  293] = -'sd2695;
    data[  294] = -'sd18865;
    data[  295] =  'sd31786;
    data[  296] =  'sd58661;
    data[  297] = -'sd80896;
    data[  298] = -'sd74749;
    data[  299] = -'sd31720;
    data[  300] = -'sd58199;
    data[  301] = -'sd79711;
    data[  302] = -'sd66454;
    data[  303] =  'sd26345;
    data[  304] =  'sd20574;
    data[  305] = -'sd19823;
    data[  306] =  'sd25080;
    data[  307] =  'sd11719;
    data[  308] = -'sd81808;
    data[  309] = -'sd81133;
    data[  310] = -'sd76408;
    data[  311] = -'sd43333;
    data[  312] =  'sd24351;
    data[  313] =  'sd6616;
    data[  314] =  'sd46312;
    data[  315] = -'sd3498;
    data[  316] = -'sd24486;
    data[  317] = -'sd7561;
    data[  318] = -'sd52927;
    data[  319] = -'sd42807;
    data[  320] =  'sd28033;
    data[  321] =  'sd32390;
    data[  322] =  'sd62889;
    data[  323] = -'sd51300;
    data[  324] = -'sd31418;
    data[  325] = -'sd56085;
    data[  326] = -'sd64913;
    data[  327] =  'sd37132;
    data[  328] = -'sd67758;
    data[  329] =  'sd17217;
    data[  330] = -'sd43322;
    data[  331] =  'sd24428;
    data[  332] =  'sd7155;
    data[  333] =  'sd50085;
    data[  334] =  'sd22913;
    data[  335] = -'sd3450;
    data[  336] = -'sd24150;
    data[  337] = -'sd5209;
    data[  338] = -'sd36463;
    data[  339] =  'sd72441;
    data[  340] =  'sd15564;
    data[  341] = -'sd54893;
    data[  342] = -'sd56569;
    data[  343] = -'sd68301;
    data[  344] =  'sd13416;
    data[  345] = -'sd69929;
    data[  346] =  'sd2020;
    data[  347] =  'sd14140;
    data[  348] = -'sd64861;
    data[  349] =  'sd37496;
    data[  350] = -'sd65210;
    data[  351] =  'sd35053;
    data[  352] =  'sd81530;
    data[  353] =  'sd79187;
    data[  354] =  'sd62786;
    data[  355] = -'sd52021;
    data[  356] = -'sd36465;
    data[  357] =  'sd72427;
    data[  358] =  'sd15466;
    data[  359] = -'sd55579;
    data[  360] = -'sd61371;
    data[  361] =  'sd61926;
    data[  362] = -'sd58041;
    data[  363] = -'sd78605;
    data[  364] = -'sd58712;
    data[  365] =  'sd80539;
    data[  366] =  'sd72250;
    data[  367] =  'sd14227;
    data[  368] = -'sd64252;
    data[  369] =  'sd41759;
    data[  370] = -'sd35369;
    data[  371] =  'sd80099;
    data[  372] =  'sd69170;
    data[  373] = -'sd7333;
    data[  374] = -'sd51331;
    data[  375] = -'sd31635;
    data[  376] = -'sd57604;
    data[  377] = -'sd75546;
    data[  378] = -'sd37299;
    data[  379] =  'sd66589;
    data[  380] = -'sd25400;
    data[  381] = -'sd13959;
    data[  382] =  'sd66128;
    data[  383] = -'sd28627;
    data[  384] = -'sd36548;
    data[  385] =  'sd71846;
    data[  386] =  'sd11399;
    data[  387] =  'sd79793;
    data[  388] =  'sd67028;
    data[  389] = -'sd22327;
    data[  390] =  'sd7552;
    data[  391] =  'sd52864;
    data[  392] =  'sd42366;
    data[  393] = -'sd31120;
    data[  394] = -'sd53999;
    data[  395] = -'sd50311;
    data[  396] = -'sd24495;
    data[  397] = -'sd7624;
    data[  398] = -'sd53368;
    data[  399] = -'sd45894;
    data[  400] =  'sd6424;
    data[  401] =  'sd44968;
    data[  402] = -'sd12906;
    data[  403] =  'sd73499;
    data[  404] =  'sd22970;
    data[  405] = -'sd3051;
    data[  406] = -'sd21357;
    data[  407] =  'sd14342;
    data[  408] = -'sd63447;
    data[  409] =  'sd47394;
    data[  410] =  'sd4076;
    data[  411] =  'sd28532;
    data[  412] =  'sd35883;
    data[  413] = -'sd76501;
    data[  414] = -'sd43984;
    data[  415] =  'sd19794;
    data[  416] = -'sd25283;
    data[  417] = -'sd13140;
    data[  418] =  'sd71861;
    data[  419] =  'sd11504;
    data[  420] =  'sd80528;
    data[  421] =  'sd72173;
    data[  422] =  'sd13688;
    data[  423] = -'sd68025;
    data[  424] =  'sd15348;
    data[  425] = -'sd56405;
    data[  426] = -'sd67153;
    data[  427] =  'sd21452;
    data[  428] = -'sd13677;
    data[  429] =  'sd68102;
    data[  430] = -'sd14809;
    data[  431] =  'sd60178;
    data[  432] = -'sd70277;
    data[  433] = -'sd416;
    data[  434] = -'sd2912;
    data[  435] = -'sd20384;
    data[  436] =  'sd21153;
    data[  437] = -'sd15770;
    data[  438] =  'sd53451;
    data[  439] =  'sd46475;
    data[  440] = -'sd2357;
    data[  441] = -'sd16499;
    data[  442] =  'sd48348;
    data[  443] =  'sd10754;
    data[  444] =  'sd75278;
    data[  445] =  'sd35423;
    data[  446] = -'sd79721;
    data[  447] = -'sd66524;
    data[  448] =  'sd25855;
    data[  449] =  'sd17144;
    data[  450] = -'sd43833;
    data[  451] =  'sd20851;
    data[  452] = -'sd17884;
    data[  453] =  'sd38653;
    data[  454] = -'sd57111;
    data[  455] = -'sd72095;
    data[  456] = -'sd13142;
    data[  457] =  'sd71847;
    data[  458] =  'sd11406;
    data[  459] =  'sd79842;
    data[  460] =  'sd67371;
    data[  461] = -'sd19926;
    data[  462] =  'sd24359;
    data[  463] =  'sd6672;
    data[  464] =  'sd46704;
    data[  465] = -'sd754;
    data[  466] = -'sd5278;
    data[  467] = -'sd36946;
    data[  468] =  'sd69060;
    data[  469] = -'sd8103;
    data[  470] = -'sd56721;
    data[  471] = -'sd69365;
    data[  472] =  'sd5968;
    data[  473] =  'sd41776;
    data[  474] = -'sd35250;
    data[  475] =  'sd80932;
    data[  476] =  'sd75001;
    data[  477] =  'sd33484;
    data[  478] =  'sd70547;
    data[  479] =  'sd2306;
    data[  480] =  'sd16142;
    data[  481] = -'sd50847;
    data[  482] = -'sd28247;
    data[  483] = -'sd33888;
    data[  484] = -'sd73375;
    data[  485] = -'sd22102;
    data[  486] =  'sd9127;
    data[  487] =  'sd63889;
    data[  488] = -'sd44300;
    data[  489] =  'sd17582;
    data[  490] = -'sd40767;
    data[  491] =  'sd42313;
    data[  492] = -'sd31491;
    data[  493] = -'sd56596;
    data[  494] = -'sd68490;
    data[  495] =  'sd12093;
    data[  496] = -'sd79190;
    data[  497] = -'sd62807;
    data[  498] =  'sd51874;
    data[  499] =  'sd35436;
    data[  500] = -'sd79630;
    data[  501] = -'sd65887;
    data[  502] =  'sd30314;
    data[  503] =  'sd48357;
    data[  504] =  'sd10817;
    data[  505] =  'sd75719;
    data[  506] =  'sd38510;
    data[  507] = -'sd58112;
    data[  508] = -'sd79102;
    data[  509] = -'sd62191;
    data[  510] =  'sd56186;
    data[  511] =  'sd65620;
    data[  512] = -'sd32183;
    data[  513] = -'sd61440;
    data[  514] =  'sd61443;
    data[  515] = -'sd61422;
    data[  516] =  'sd61569;
    data[  517] = -'sd60540;
    data[  518] =  'sd67743;
    data[  519] = -'sd17322;
    data[  520] =  'sd42587;
    data[  521] = -'sd29573;
    data[  522] = -'sd43170;
    data[  523] =  'sd25492;
    data[  524] =  'sd14603;
    data[  525] = -'sd61620;
    data[  526] =  'sd60183;
    data[  527] = -'sd70242;
    data[  528] = -'sd171;
    data[  529] = -'sd1197;
    data[  530] = -'sd8379;
    data[  531] = -'sd58653;
    data[  532] =  'sd80952;
    data[  533] =  'sd75141;
    data[  534] =  'sd34464;
    data[  535] =  'sd77407;
    data[  536] =  'sd50326;
    data[  537] =  'sd24600;
    data[  538] =  'sd8359;
    data[  539] =  'sd58513;
    data[  540] =  'sd81909;
    data[  541] =  'sd81840;
    data[  542] =  'sd81357;
    data[  543] =  'sd77976;
    data[  544] =  'sd54309;
    data[  545] =  'sd52481;
    data[  546] =  'sd39685;
    data[  547] = -'sd49887;
    data[  548] = -'sd21527;
    data[  549] =  'sd13152;
    data[  550] = -'sd71777;
    data[  551] = -'sd10916;
    data[  552] = -'sd76412;
    data[  553] = -'sd43361;
    data[  554] =  'sd24155;
    data[  555] =  'sd5244;
    data[  556] =  'sd36708;
    data[  557] = -'sd70726;
    data[  558] = -'sd3559;
    data[  559] = -'sd24913;
    data[  560] = -'sd10550;
    data[  561] = -'sd73850;
    data[  562] = -'sd25427;
    data[  563] = -'sd14148;
    data[  564] =  'sd64805;
    data[  565] = -'sd37888;
    data[  566] =  'sd62466;
    data[  567] = -'sd54261;
    data[  568] = -'sd52145;
    data[  569] = -'sd37333;
    data[  570] =  'sd66351;
    data[  571] = -'sd27066;
    data[  572] = -'sd25621;
    data[  573] = -'sd15506;
    data[  574] =  'sd55299;
    data[  575] =  'sd59411;
    data[  576] = -'sd75646;
    data[  577] = -'sd37999;
    data[  578] =  'sd61689;
    data[  579] = -'sd59700;
    data[  580] =  'sd73623;
    data[  581] =  'sd23838;
    data[  582] =  'sd3025;
    data[  583] =  'sd21175;
    data[  584] = -'sd15616;
    data[  585] =  'sd54529;
    data[  586] =  'sd54021;
    data[  587] =  'sd50465;
    data[  588] =  'sd25573;
    data[  589] =  'sd15170;
    data[  590] = -'sd57651;
    data[  591] = -'sd75875;
    data[  592] = -'sd39602;
    data[  593] =  'sd50468;
    data[  594] =  'sd25594;
    data[  595] =  'sd15317;
    data[  596] = -'sd56622;
    data[  597] = -'sd68672;
    data[  598] =  'sd10819;
    data[  599] =  'sd75733;
    data[  600] =  'sd38608;
    data[  601] = -'sd57426;
    data[  602] = -'sd74300;
    data[  603] = -'sd28577;
    data[  604] = -'sd36198;
    data[  605] =  'sd74296;
    data[  606] =  'sd28549;
    data[  607] =  'sd36002;
    data[  608] = -'sd75668;
    data[  609] = -'sd38153;
    data[  610] =  'sd60611;
    data[  611] = -'sd67246;
    data[  612] =  'sd20801;
    data[  613] = -'sd18234;
    data[  614] =  'sd36203;
    data[  615] = -'sd74261;
    data[  616] = -'sd28304;
    data[  617] = -'sd34287;
    data[  618] = -'sd76168;
    data[  619] = -'sd41653;
    data[  620] =  'sd36111;
    data[  621] = -'sd74905;
    data[  622] = -'sd32812;
    data[  623] = -'sd65843;
    data[  624] =  'sd30622;
    data[  625] =  'sd50513;
    data[  626] =  'sd25909;
    data[  627] =  'sd17522;
    data[  628] = -'sd41187;
    data[  629] =  'sd39373;
    data[  630] = -'sd52071;
    data[  631] = -'sd36815;
    data[  632] =  'sd69977;
    data[  633] = -'sd1684;
    data[  634] = -'sd11788;
    data[  635] =  'sd81325;
    data[  636] =  'sd77752;
    data[  637] =  'sd52741;
    data[  638] =  'sd41505;
    data[  639] = -'sd37147;
    data[  640] =  'sd67653;
    data[  641] = -'sd17952;
    data[  642] =  'sd38177;
    data[  643] = -'sd60443;
    data[  644] =  'sd68422;
    data[  645] = -'sd12569;
    data[  646] =  'sd75858;
    data[  647] =  'sd39483;
    data[  648] = -'sd51301;
    data[  649] = -'sd31425;
    data[  650] = -'sd56134;
    data[  651] = -'sd65256;
    data[  652] =  'sd34731;
    data[  653] =  'sd79276;
    data[  654] =  'sd63409;
    data[  655] = -'sd47660;
    data[  656] = -'sd5938;
    data[  657] = -'sd41566;
    data[  658] =  'sd36720;
    data[  659] = -'sd70642;
    data[  660] = -'sd2971;
    data[  661] = -'sd20797;
    data[  662] =  'sd18262;
    data[  663] = -'sd36007;
    data[  664] =  'sd75633;
    data[  665] =  'sd37908;
    data[  666] = -'sd62326;
    data[  667] =  'sd55241;
    data[  668] =  'sd59005;
    data[  669] = -'sd78488;
    data[  670] = -'sd57893;
    data[  671] = -'sd77569;
    data[  672] = -'sd51460;
    data[  673] = -'sd32538;
    data[  674] = -'sd63925;
    data[  675] =  'sd44048;
    data[  676] = -'sd19346;
    data[  677] =  'sd28419;
    data[  678] =  'sd35092;
    data[  679] =  'sd81803;
    data[  680] =  'sd81098;
    data[  681] =  'sd76163;
    data[  682] =  'sd41618;
    data[  683] = -'sd36356;
    data[  684] =  'sd73190;
    data[  685] =  'sd20807;
    data[  686] = -'sd18192;
    data[  687] =  'sd36497;
    data[  688] = -'sd72203;
    data[  689] = -'sd13898;
    data[  690] =  'sd66555;
    data[  691] = -'sd25638;
    data[  692] = -'sd15625;
    data[  693] =  'sd54466;
    data[  694] =  'sd53580;
    data[  695] =  'sd47378;
    data[  696] =  'sd3964;
    data[  697] =  'sd27748;
    data[  698] =  'sd30395;
    data[  699] =  'sd48924;
    data[  700] =  'sd14786;
    data[  701] = -'sd60339;
    data[  702] =  'sd69150;
    data[  703] = -'sd7473;
    data[  704] = -'sd52311;
    data[  705] = -'sd38495;
    data[  706] =  'sd58217;
    data[  707] =  'sd79837;
    data[  708] =  'sd67336;
    data[  709] = -'sd20171;
    data[  710] =  'sd22644;
    data[  711] = -'sd5333;
    data[  712] = -'sd37331;
    data[  713] =  'sd66365;
    data[  714] = -'sd26968;
    data[  715] = -'sd24935;
    data[  716] = -'sd10704;
    data[  717] = -'sd74928;
    data[  718] = -'sd32973;
    data[  719] = -'sd66970;
    data[  720] =  'sd22733;
    data[  721] = -'sd4710;
    data[  722] = -'sd32970;
    data[  723] = -'sd66949;
    data[  724] =  'sd22880;
    data[  725] = -'sd3681;
    data[  726] = -'sd25767;
    data[  727] = -'sd16528;
    data[  728] =  'sd48145;
    data[  729] =  'sd9333;
    data[  730] =  'sd65331;
    data[  731] = -'sd34206;
    data[  732] = -'sd75601;
    data[  733] = -'sd37684;
    data[  734] =  'sd63894;
    data[  735] = -'sd44265;
    data[  736] =  'sd17827;
    data[  737] = -'sd39052;
    data[  738] =  'sd54318;
    data[  739] =  'sd52544;
    data[  740] =  'sd40126;
    data[  741] = -'sd46800;
    data[  742] =  'sd82;
    data[  743] =  'sd574;
    data[  744] =  'sd4018;
    data[  745] =  'sd28126;
    data[  746] =  'sd33041;
    data[  747] =  'sd67446;
    data[  748] = -'sd19401;
    data[  749] =  'sd28034;
    data[  750] =  'sd32397;
    data[  751] =  'sd62938;
    data[  752] = -'sd50957;
    data[  753] = -'sd29017;
    data[  754] = -'sd39278;
    data[  755] =  'sd52736;
    data[  756] =  'sd41470;
    data[  757] = -'sd37392;
    data[  758] =  'sd65938;
    data[  759] = -'sd29957;
    data[  760] = -'sd45858;
    data[  761] =  'sd6676;
    data[  762] =  'sd46732;
    data[  763] = -'sd558;
    data[  764] = -'sd3906;
    data[  765] = -'sd27342;
    data[  766] = -'sd27553;
    data[  767] = -'sd29030;
    data[  768] = -'sd39369;
    data[  769] =  'sd52099;
    data[  770] =  'sd37011;
    data[  771] = -'sd68605;
    data[  772] =  'sd11288;
    data[  773] =  'sd79016;
    data[  774] =  'sd61589;
    data[  775] = -'sd60400;
    data[  776] =  'sd68723;
    data[  777] = -'sd10462;
    data[  778] = -'sd73234;
    data[  779] = -'sd21115;
    data[  780] =  'sd16036;
    data[  781] = -'sd51589;
    data[  782] = -'sd33441;
    data[  783] = -'sd70246;
    data[  784] = -'sd199;
    data[  785] = -'sd1393;
    data[  786] = -'sd9751;
    data[  787] = -'sd68257;
    data[  788] =  'sd13724;
    data[  789] = -'sd67773;
    data[  790] =  'sd17112;
    data[  791] = -'sd44057;
    data[  792] =  'sd19283;
    data[  793] = -'sd28860;
    data[  794] = -'sd38179;
    data[  795] =  'sd60429;
    data[  796] = -'sd68520;
    data[  797] =  'sd11883;
    data[  798] = -'sd80660;
    data[  799] = -'sd73097;
    data[  800] = -'sd20156;
    data[  801] =  'sd22749;
    data[  802] = -'sd4598;
    data[  803] = -'sd32186;
    data[  804] = -'sd61461;
    data[  805] =  'sd61296;
    data[  806] = -'sd62451;
    data[  807] =  'sd54366;
    data[  808] =  'sd52880;
    data[  809] =  'sd42478;
    data[  810] = -'sd30336;
    data[  811] = -'sd48511;
    data[  812] = -'sd11895;
    data[  813] =  'sd80576;
    data[  814] =  'sd72509;
    data[  815] =  'sd16040;
    data[  816] = -'sd51561;
    data[  817] = -'sd33245;
    data[  818] = -'sd68874;
    data[  819] =  'sd9405;
    data[  820] =  'sd65835;
    data[  821] = -'sd30678;
    data[  822] = -'sd50905;
    data[  823] = -'sd28653;
    data[  824] = -'sd36730;
    data[  825] =  'sd70572;
    data[  826] =  'sd2481;
    data[  827] =  'sd17367;
    data[  828] = -'sd42272;
    data[  829] =  'sd31778;
    data[  830] =  'sd58605;
    data[  831] = -'sd81288;
    data[  832] = -'sd77493;
    data[  833] = -'sd50928;
    data[  834] = -'sd28814;
    data[  835] = -'sd37857;
    data[  836] =  'sd62683;
    data[  837] = -'sd52742;
    data[  838] = -'sd41512;
    data[  839] =  'sd37098;
    data[  840] = -'sd67996;
    data[  841] =  'sd15551;
    data[  842] = -'sd54984;
    data[  843] = -'sd57206;
    data[  844] = -'sd72760;
    data[  845] = -'sd17797;
    data[  846] =  'sd39262;
    data[  847] = -'sd52848;
    data[  848] = -'sd42254;
    data[  849] =  'sd31904;
    data[  850] =  'sd59487;
    data[  851] = -'sd75114;
    data[  852] = -'sd34275;
    data[  853] = -'sd76084;
    data[  854] = -'sd41065;
    data[  855] =  'sd40227;
    data[  856] = -'sd46093;
    data[  857] =  'sd5031;
    data[  858] =  'sd35217;
    data[  859] = -'sd81163;
    data[  860] = -'sd76618;
    data[  861] = -'sd44803;
    data[  862] =  'sd14061;
    data[  863] = -'sd65414;
    data[  864] =  'sd33625;
    data[  865] =  'sd71534;
    data[  866] =  'sd9215;
    data[  867] =  'sd64505;
    data[  868] = -'sd39988;
    data[  869] =  'sd47766;
    data[  870] =  'sd6680;
    data[  871] =  'sd46760;
    data[  872] = -'sd362;
    data[  873] = -'sd2534;
    data[  874] = -'sd17738;
    data[  875] =  'sd39675;
    data[  876] = -'sd49957;
    data[  877] = -'sd22017;
    data[  878] =  'sd9722;
    data[  879] =  'sd68054;
    data[  880] = -'sd15145;
    data[  881] =  'sd57826;
    data[  882] =  'sd77100;
    data[  883] =  'sd48177;
    data[  884] =  'sd9557;
    data[  885] =  'sd66899;
    data[  886] = -'sd23230;
    data[  887] =  'sd1231;
    data[  888] =  'sd8617;
    data[  889] =  'sd60319;
    data[  890] = -'sd69290;
    data[  891] =  'sd6493;
    data[  892] =  'sd45451;
    data[  893] = -'sd9525;
    data[  894] = -'sd66675;
    data[  895] =  'sd24798;
    data[  896] =  'sd9745;
    data[  897] =  'sd68215;
    data[  898] = -'sd14018;
    data[  899] =  'sd65715;
    data[  900] = -'sd31518;
    data[  901] = -'sd56785;
    data[  902] = -'sd69813;
    data[  903] =  'sd2832;
    data[  904] =  'sd19824;
    data[  905] = -'sd25073;
    data[  906] = -'sd11670;
    data[  907] = -'sd81690;
    data[  908] = -'sd80307;
    data[  909] = -'sd70626;
    data[  910] = -'sd2859;
    data[  911] = -'sd20013;
    data[  912] =  'sd23750;
    data[  913] =  'sd2409;
    data[  914] =  'sd16863;
    data[  915] = -'sd45800;
    data[  916] =  'sd7082;
    data[  917] =  'sd49574;
    data[  918] =  'sd19336;
    data[  919] = -'sd28489;
    data[  920] = -'sd35582;
    data[  921] =  'sd78608;
    data[  922] =  'sd58733;
    data[  923] = -'sd80392;
    data[  924] = -'sd71221;
    data[  925] = -'sd7024;
    data[  926] = -'sd49168;
    data[  927] = -'sd16494;
    data[  928] =  'sd48383;
    data[  929] =  'sd10999;
    data[  930] =  'sd76993;
    data[  931] =  'sd47428;
    data[  932] =  'sd4314;
    data[  933] =  'sd30198;
    data[  934] =  'sd47545;
    data[  935] =  'sd5133;
    data[  936] =  'sd35931;
    data[  937] = -'sd76165;
    data[  938] = -'sd41632;
    data[  939] =  'sd36258;
    data[  940] = -'sd73876;
    data[  941] = -'sd25609;
    data[  942] = -'sd15422;
    data[  943] =  'sd55887;
    data[  944] =  'sd63527;
    data[  945] = -'sd46834;
    data[  946] = -'sd156;
    data[  947] = -'sd1092;
    data[  948] = -'sd7644;
    data[  949] = -'sd53508;
    data[  950] = -'sd46874;
    data[  951] = -'sd436;
    data[  952] = -'sd3052;
    data[  953] = -'sd21364;
    data[  954] =  'sd14293;
    data[  955] = -'sd63790;
    data[  956] =  'sd44993;
    data[  957] = -'sd12731;
    data[  958] =  'sd74724;
    data[  959] =  'sd31545;
    data[  960] =  'sd56974;
    data[  961] =  'sd71136;
    data[  962] =  'sd6429;
    data[  963] =  'sd45003;
    data[  964] = -'sd12661;
    data[  965] =  'sd75214;
    data[  966] =  'sd34975;
    data[  967] =  'sd80984;
    data[  968] =  'sd75365;
    data[  969] =  'sd36032;
    data[  970] = -'sd75458;
    data[  971] = -'sd36683;
    data[  972] =  'sd70901;
    data[  973] =  'sd4784;
    data[  974] =  'sd33488;
    data[  975] =  'sd70575;
    data[  976] =  'sd2502;
    data[  977] =  'sd17514;
    data[  978] = -'sd41243;
    data[  979] =  'sd38981;
    data[  980] = -'sd54815;
    data[  981] = -'sd56023;
    data[  982] = -'sd64479;
    data[  983] =  'sd40170;
    data[  984] = -'sd46492;
    data[  985] =  'sd2238;
    data[  986] =  'sd15666;
    data[  987] = -'sd54179;
    data[  988] = -'sd51571;
    data[  989] = -'sd33315;
    data[  990] = -'sd69364;
    data[  991] =  'sd5975;
    data[  992] =  'sd41825;
    data[  993] = -'sd34907;
    data[  994] = -'sd80508;
    data[  995] = -'sd72033;
    data[  996] = -'sd12708;
    data[  997] =  'sd74885;
    data[  998] =  'sd32672;
    data[  999] =  'sd64863;
    data[ 1000] = -'sd37482;
    data[ 1001] =  'sd65308;
    data[ 1002] = -'sd34367;
    data[ 1003] = -'sd76728;
    data[ 1004] = -'sd45573;
    data[ 1005] =  'sd8671;
    data[ 1006] =  'sd60697;
    data[ 1007] = -'sd66644;
    data[ 1008] =  'sd25015;
    data[ 1009] =  'sd11264;
    data[ 1010] =  'sd78848;
    data[ 1011] =  'sd60413;
    data[ 1012] = -'sd68632;
    data[ 1013] =  'sd11099;
    data[ 1014] =  'sd77693;
    data[ 1015] =  'sd52328;
    data[ 1016] =  'sd38614;
    data[ 1017] = -'sd57384;
    data[ 1018] = -'sd74006;
    data[ 1019] = -'sd26519;
    data[ 1020] = -'sd21792;
    data[ 1021] =  'sd11297;
    data[ 1022] =  'sd79079;
    data[ 1023] =  'sd62030;
    data[ 1024] = -'sd57313;
    data[ 1025] = -'sd73509;
    data[ 1026] = -'sd23040;
    data[ 1027] =  'sd2561;
    data[ 1028] =  'sd17927;
    data[ 1029] = -'sd38352;
    data[ 1030] =  'sd59218;
    data[ 1031] = -'sd76997;
    data[ 1032] = -'sd47456;
    data[ 1033] = -'sd4510;
    data[ 1034] = -'sd31570;
    data[ 1035] = -'sd57149;
    data[ 1036] = -'sd72361;
    data[ 1037] = -'sd15004;
    data[ 1038] =  'sd58813;
    data[ 1039] = -'sd79832;
    data[ 1040] = -'sd67301;
    data[ 1041] =  'sd20416;
    data[ 1042] = -'sd20929;
    data[ 1043] =  'sd17338;
    data[ 1044] = -'sd42475;
    data[ 1045] =  'sd30357;
    data[ 1046] =  'sd48658;
    data[ 1047] =  'sd12924;
    data[ 1048] = -'sd73373;
    data[ 1049] = -'sd22088;
    data[ 1050] =  'sd9225;
    data[ 1051] =  'sd64575;
    data[ 1052] = -'sd39498;
    data[ 1053] =  'sd51196;
    data[ 1054] =  'sd30690;
    data[ 1055] =  'sd50989;
    data[ 1056] =  'sd29241;
    data[ 1057] =  'sd40846;
    data[ 1058] = -'sd41760;
    data[ 1059] =  'sd35362;
    data[ 1060] = -'sd80148;
    data[ 1061] = -'sd69513;
    data[ 1062] =  'sd4932;
    data[ 1063] =  'sd34524;
    data[ 1064] =  'sd77827;
    data[ 1065] =  'sd53266;
    data[ 1066] =  'sd45180;
    data[ 1067] = -'sd11422;
    data[ 1068] = -'sd79954;
    data[ 1069] = -'sd68155;
    data[ 1070] =  'sd14438;
    data[ 1071] = -'sd62775;
    data[ 1072] =  'sd52098;
    data[ 1073] =  'sd37004;
    data[ 1074] = -'sd68654;
    data[ 1075] =  'sd10945;
    data[ 1076] =  'sd76615;
    data[ 1077] =  'sd44782;
    data[ 1078] = -'sd14208;
    data[ 1079] =  'sd64385;
    data[ 1080] = -'sd40828;
    data[ 1081] =  'sd41886;
    data[ 1082] = -'sd34480;
    data[ 1083] = -'sd77519;
    data[ 1084] = -'sd51110;
    data[ 1085] = -'sd30088;
    data[ 1086] = -'sd46775;
    data[ 1087] =  'sd257;
    data[ 1088] =  'sd1799;
    data[ 1089] =  'sd12593;
    data[ 1090] = -'sd75690;
    data[ 1091] = -'sd38307;
    data[ 1092] =  'sd59533;
    data[ 1093] = -'sd74792;
    data[ 1094] = -'sd32021;
    data[ 1095] = -'sd60306;
    data[ 1096] =  'sd69381;
    data[ 1097] = -'sd5856;
    data[ 1098] = -'sd40992;
    data[ 1099] =  'sd40738;
    data[ 1100] = -'sd42516;
    data[ 1101] =  'sd30070;
    data[ 1102] =  'sd46649;
    data[ 1103] = -'sd1139;
    data[ 1104] = -'sd7973;
    data[ 1105] = -'sd55811;
    data[ 1106] = -'sd62995;
    data[ 1107] =  'sd50558;
    data[ 1108] =  'sd26224;
    data[ 1109] =  'sd19727;
    data[ 1110] = -'sd25752;
    data[ 1111] = -'sd16423;
    data[ 1112] =  'sd48880;
    data[ 1113] =  'sd14478;
    data[ 1114] = -'sd62495;
    data[ 1115] =  'sd54058;
    data[ 1116] =  'sd50724;
    data[ 1117] =  'sd27386;
    data[ 1118] =  'sd27861;
    data[ 1119] =  'sd31186;
    data[ 1120] =  'sd54461;
    data[ 1121] =  'sd53545;
    data[ 1122] =  'sd47133;
    data[ 1123] =  'sd2249;
    data[ 1124] =  'sd15743;
    data[ 1125] = -'sd53640;
    data[ 1126] = -'sd47798;
    data[ 1127] = -'sd6904;
    data[ 1128] = -'sd48328;
    data[ 1129] = -'sd10614;
    data[ 1130] = -'sd74298;
    data[ 1131] = -'sd28563;
    data[ 1132] = -'sd36100;
    data[ 1133] =  'sd74982;
    data[ 1134] =  'sd33351;
    data[ 1135] =  'sd69616;
    data[ 1136] = -'sd4211;
    data[ 1137] = -'sd29477;
    data[ 1138] = -'sd42498;
    data[ 1139] =  'sd30196;
    data[ 1140] =  'sd47531;
    data[ 1141] =  'sd5035;
    data[ 1142] =  'sd35245;
    data[ 1143] = -'sd80967;
    data[ 1144] = -'sd75246;
    data[ 1145] = -'sd35199;
    data[ 1146] =  'sd81289;
    data[ 1147] =  'sd77500;
    data[ 1148] =  'sd50977;
    data[ 1149] =  'sd29157;
    data[ 1150] =  'sd40258;
    data[ 1151] = -'sd45876;
    data[ 1152] =  'sd6550;
    data[ 1153] =  'sd45850;
    data[ 1154] = -'sd6732;
    data[ 1155] = -'sd47124;
    data[ 1156] = -'sd2186;
    data[ 1157] = -'sd15302;
    data[ 1158] =  'sd56727;
    data[ 1159] =  'sd69407;
    data[ 1160] = -'sd5674;
    data[ 1161] = -'sd39718;
    data[ 1162] =  'sd49656;
    data[ 1163] =  'sd19910;
    data[ 1164] = -'sd24471;
    data[ 1165] = -'sd7456;
    data[ 1166] = -'sd52192;
    data[ 1167] = -'sd37662;
    data[ 1168] =  'sd64048;
    data[ 1169] = -'sd43187;
    data[ 1170] =  'sd25373;
    data[ 1171] =  'sd13770;
    data[ 1172] = -'sd67451;
    data[ 1173] =  'sd19366;
    data[ 1174] = -'sd28279;
    data[ 1175] = -'sd34112;
    data[ 1176] = -'sd74943;
    data[ 1177] = -'sd33078;
    data[ 1178] = -'sd67705;
    data[ 1179] =  'sd17588;
    data[ 1180] = -'sd40725;
    data[ 1181] =  'sd42607;
    data[ 1182] = -'sd29433;
    data[ 1183] = -'sd42190;
    data[ 1184] =  'sd32352;
    data[ 1185] =  'sd62623;
    data[ 1186] = -'sd53162;
    data[ 1187] = -'sd44452;
    data[ 1188] =  'sd16518;
    data[ 1189] = -'sd48215;
    data[ 1190] = -'sd9823;
    data[ 1191] = -'sd68761;
    data[ 1192] =  'sd10196;
    data[ 1193] =  'sd71372;
    data[ 1194] =  'sd8081;
    data[ 1195] =  'sd56567;
    data[ 1196] =  'sd68287;
    data[ 1197] = -'sd13514;
    data[ 1198] =  'sd69243;
    data[ 1199] = -'sd6822;
    data[ 1200] = -'sd47754;
    data[ 1201] = -'sd6596;
    data[ 1202] = -'sd46172;
    data[ 1203] =  'sd4478;
    data[ 1204] =  'sd31346;
    data[ 1205] =  'sd55581;
    data[ 1206] =  'sd61385;
    data[ 1207] = -'sd61828;
    data[ 1208] =  'sd58727;
    data[ 1209] = -'sd80434;
    data[ 1210] = -'sd71515;
    data[ 1211] = -'sd9082;
    data[ 1212] = -'sd63574;
    data[ 1213] =  'sd46505;
    data[ 1214] = -'sd2147;
    data[ 1215] = -'sd15029;
    data[ 1216] =  'sd58638;
    data[ 1217] = -'sd81057;
    data[ 1218] = -'sd75876;
    data[ 1219] = -'sd39609;
    data[ 1220] =  'sd50419;
    data[ 1221] =  'sd25251;
    data[ 1222] =  'sd12916;
    data[ 1223] = -'sd73429;
    data[ 1224] = -'sd22480;
    data[ 1225] =  'sd6481;
    data[ 1226] =  'sd45367;
    data[ 1227] = -'sd10113;
    data[ 1228] = -'sd70791;
    data[ 1229] = -'sd4014;
    data[ 1230] = -'sd28098;
    data[ 1231] = -'sd32845;
    data[ 1232] = -'sd66074;
    data[ 1233] =  'sd29005;
    data[ 1234] =  'sd39194;
    data[ 1235] = -'sd53324;
    data[ 1236] = -'sd45586;
    data[ 1237] =  'sd8580;
    data[ 1238] =  'sd60060;
    data[ 1239] = -'sd71103;
    data[ 1240] = -'sd6198;
    data[ 1241] = -'sd43386;
    data[ 1242] =  'sd23980;
    data[ 1243] =  'sd4019;
    data[ 1244] =  'sd28133;
    data[ 1245] =  'sd33090;
    data[ 1246] =  'sd67789;
    data[ 1247] = -'sd17000;
    data[ 1248] =  'sd44841;
    data[ 1249] = -'sd13795;
    data[ 1250] =  'sd67276;
    data[ 1251] = -'sd20591;
    data[ 1252] =  'sd19704;
    data[ 1253] = -'sd25913;
    data[ 1254] = -'sd17550;
    data[ 1255] =  'sd40991;
    data[ 1256] = -'sd40745;
    data[ 1257] =  'sd42467;
    data[ 1258] = -'sd30413;
    data[ 1259] = -'sd49050;
    data[ 1260] = -'sd15668;
    data[ 1261] =  'sd54165;
    data[ 1262] =  'sd51473;
    data[ 1263] =  'sd32629;
    data[ 1264] =  'sd64562;
    data[ 1265] = -'sd39589;
    data[ 1266] =  'sd50559;
    data[ 1267] =  'sd26231;
    data[ 1268] =  'sd19776;
    data[ 1269] = -'sd25409;
    data[ 1270] = -'sd14022;
    data[ 1271] =  'sd65687;
    data[ 1272] = -'sd31714;
    data[ 1273] = -'sd58157;
    data[ 1274] = -'sd79417;
    data[ 1275] = -'sd64396;
    data[ 1276] =  'sd40751;
    data[ 1277] = -'sd42425;
    data[ 1278] =  'sd30707;
    data[ 1279] =  'sd51108;
    data[ 1280] =  'sd30074;
    data[ 1281] =  'sd46677;
    data[ 1282] = -'sd943;
    data[ 1283] = -'sd6601;
    data[ 1284] = -'sd46207;
    data[ 1285] =  'sd4233;
    data[ 1286] =  'sd29631;
    data[ 1287] =  'sd43576;
    data[ 1288] = -'sd22650;
    data[ 1289] =  'sd5291;
    data[ 1290] =  'sd37037;
    data[ 1291] = -'sd68423;
    data[ 1292] =  'sd12562;
    data[ 1293] = -'sd75907;
    data[ 1294] = -'sd39826;
    data[ 1295] =  'sd48900;
    data[ 1296] =  'sd14618;
    data[ 1297] = -'sd61515;
    data[ 1298] =  'sd60918;
    data[ 1299] = -'sd65097;
    data[ 1300] =  'sd35844;
    data[ 1301] = -'sd76774;
    data[ 1302] = -'sd45895;
    data[ 1303] =  'sd6417;
    data[ 1304] =  'sd44919;
    data[ 1305] = -'sd13249;
    data[ 1306] =  'sd71098;
    data[ 1307] =  'sd6163;
    data[ 1308] =  'sd43141;
    data[ 1309] = -'sd25695;
    data[ 1310] = -'sd16024;
    data[ 1311] =  'sd51673;
    data[ 1312] =  'sd34029;
    data[ 1313] =  'sd74362;
    data[ 1314] =  'sd29011;
    data[ 1315] =  'sd39236;
    data[ 1316] = -'sd53030;
    data[ 1317] = -'sd43528;
    data[ 1318] =  'sd22986;
    data[ 1319] = -'sd2939;
    data[ 1320] = -'sd20573;
    data[ 1321] =  'sd19830;
    data[ 1322] = -'sd25031;
    data[ 1323] = -'sd11376;
    data[ 1324] = -'sd79632;
    data[ 1325] = -'sd65901;
    data[ 1326] =  'sd30216;
    data[ 1327] =  'sd47671;
    data[ 1328] =  'sd6015;
    data[ 1329] =  'sd42105;
    data[ 1330] = -'sd32947;
    data[ 1331] = -'sd66788;
    data[ 1332] =  'sd24007;
    data[ 1333] =  'sd4208;
    data[ 1334] =  'sd29456;
    data[ 1335] =  'sd42351;
    data[ 1336] = -'sd31225;
    data[ 1337] = -'sd54734;
    data[ 1338] = -'sd55456;
    data[ 1339] = -'sd60510;
    data[ 1340] =  'sd67953;
    data[ 1341] = -'sd15852;
    data[ 1342] =  'sd52877;
    data[ 1343] =  'sd42457;
    data[ 1344] = -'sd30483;
    data[ 1345] = -'sd49540;
    data[ 1346] = -'sd19098;
    data[ 1347] =  'sd30155;
    data[ 1348] =  'sd47244;
    data[ 1349] =  'sd3026;
    data[ 1350] =  'sd21182;
    data[ 1351] = -'sd15567;
    data[ 1352] =  'sd54872;
    data[ 1353] =  'sd56422;
    data[ 1354] =  'sd67272;
    data[ 1355] = -'sd20619;
    data[ 1356] =  'sd19508;
    data[ 1357] = -'sd27285;
    data[ 1358] = -'sd27154;
    data[ 1359] = -'sd26237;
    data[ 1360] = -'sd19818;
    data[ 1361] =  'sd25115;
    data[ 1362] =  'sd11964;
    data[ 1363] = -'sd80093;
    data[ 1364] = -'sd69128;
    data[ 1365] =  'sd7627;
    data[ 1366] =  'sd53389;
    data[ 1367] =  'sd46041;
    data[ 1368] = -'sd5395;
    data[ 1369] = -'sd37765;
    data[ 1370] =  'sd63327;
    data[ 1371] = -'sd48234;
    data[ 1372] = -'sd9956;
    data[ 1373] = -'sd69692;
    data[ 1374] =  'sd3679;
    data[ 1375] =  'sd25753;
    data[ 1376] =  'sd16430;
    data[ 1377] = -'sd48831;
    data[ 1378] = -'sd14135;
    data[ 1379] =  'sd64896;
    data[ 1380] = -'sd37251;
    data[ 1381] =  'sd66925;
    data[ 1382] = -'sd23048;
    data[ 1383] =  'sd2505;
    data[ 1384] =  'sd17535;
    data[ 1385] = -'sd41096;
    data[ 1386] =  'sd40010;
    data[ 1387] = -'sd47612;
    data[ 1388] = -'sd5602;
    data[ 1389] = -'sd39214;
    data[ 1390] =  'sd53184;
    data[ 1391] =  'sd44606;
    data[ 1392] = -'sd15440;
    data[ 1393] =  'sd55761;
    data[ 1394] =  'sd62645;
    data[ 1395] = -'sd53008;
    data[ 1396] = -'sd43374;
    data[ 1397] =  'sd24064;
    data[ 1398] =  'sd4607;
    data[ 1399] =  'sd32249;
    data[ 1400] =  'sd61902;
    data[ 1401] = -'sd58209;
    data[ 1402] = -'sd79781;
    data[ 1403] = -'sd66944;
    data[ 1404] =  'sd22915;
    data[ 1405] = -'sd3436;
    data[ 1406] = -'sd24052;
    data[ 1407] = -'sd4523;
    data[ 1408] = -'sd31661;
    data[ 1409] = -'sd57786;
    data[ 1410] = -'sd76820;
    data[ 1411] = -'sd46217;
    data[ 1412] =  'sd4163;
    data[ 1413] =  'sd29141;
    data[ 1414] =  'sd40146;
    data[ 1415] = -'sd46660;
    data[ 1416] =  'sd1062;
    data[ 1417] =  'sd7434;
    data[ 1418] =  'sd52038;
    data[ 1419] =  'sd36584;
    data[ 1420] = -'sd71594;
    data[ 1421] = -'sd9635;
    data[ 1422] = -'sd67445;
    data[ 1423] =  'sd19408;
    data[ 1424] = -'sd27985;
    data[ 1425] = -'sd32054;
    data[ 1426] = -'sd60537;
    data[ 1427] =  'sd67764;
    data[ 1428] = -'sd17175;
    data[ 1429] =  'sd43616;
    data[ 1430] = -'sd22370;
    data[ 1431] =  'sd7251;
    data[ 1432] =  'sd50757;
    data[ 1433] =  'sd27617;
    data[ 1434] =  'sd29478;
    data[ 1435] =  'sd42505;
    data[ 1436] = -'sd30147;
    data[ 1437] = -'sd47188;
    data[ 1438] = -'sd2634;
    data[ 1439] = -'sd18438;
    data[ 1440] =  'sd34775;
    data[ 1441] =  'sd79584;
    data[ 1442] =  'sd65565;
    data[ 1443] = -'sd32568;
    data[ 1444] = -'sd64135;
    data[ 1445] =  'sd42578;
    data[ 1446] = -'sd29636;
    data[ 1447] = -'sd43611;
    data[ 1448] =  'sd22405;
    data[ 1449] = -'sd7006;
    data[ 1450] = -'sd49042;
    data[ 1451] = -'sd15612;
    data[ 1452] =  'sd54557;
    data[ 1453] =  'sd54217;
    data[ 1454] =  'sd51837;
    data[ 1455] =  'sd35177;
    data[ 1456] = -'sd81443;
    data[ 1457] = -'sd78578;
    data[ 1458] = -'sd58523;
    data[ 1459] =  'sd81862;
    data[ 1460] =  'sd81511;
    data[ 1461] =  'sd79054;
    data[ 1462] =  'sd61855;
    data[ 1463] = -'sd58538;
    data[ 1464] =  'sd81757;
    data[ 1465] =  'sd80776;
    data[ 1466] =  'sd73909;
    data[ 1467] =  'sd25840;
    data[ 1468] =  'sd17039;
    data[ 1469] = -'sd44568;
    data[ 1470] =  'sd15706;
    data[ 1471] = -'sd53899;
    data[ 1472] = -'sd49611;
    data[ 1473] = -'sd19595;
    data[ 1474] =  'sd26676;
    data[ 1475] =  'sd22891;
    data[ 1476] = -'sd3604;
    data[ 1477] = -'sd25228;
    data[ 1478] = -'sd12755;
    data[ 1479] =  'sd74556;
    data[ 1480] =  'sd30369;
    data[ 1481] =  'sd48742;
    data[ 1482] =  'sd13512;
    data[ 1483] = -'sd69257;
    data[ 1484] =  'sd6724;
    data[ 1485] =  'sd47068;
    data[ 1486] =  'sd1794;
    data[ 1487] =  'sd12558;
    data[ 1488] = -'sd75935;
    data[ 1489] = -'sd40022;
    data[ 1490] =  'sd47528;
    data[ 1491] =  'sd5014;
    data[ 1492] =  'sd35098;
    data[ 1493] =  'sd81845;
    data[ 1494] =  'sd81392;
    data[ 1495] =  'sd78221;
    data[ 1496] =  'sd56024;
    data[ 1497] =  'sd64486;
    data[ 1498] = -'sd40121;
    data[ 1499] =  'sd46835;
    data[ 1500] =  'sd163;
    data[ 1501] =  'sd1141;
    data[ 1502] =  'sd7987;
    data[ 1503] =  'sd55909;
    data[ 1504] =  'sd63681;
    data[ 1505] = -'sd45756;
    data[ 1506] =  'sd7390;
    data[ 1507] =  'sd51730;
    data[ 1508] =  'sd34428;
    data[ 1509] =  'sd77155;
    data[ 1510] =  'sd48562;
    data[ 1511] =  'sd12252;
    data[ 1512] = -'sd78077;
    data[ 1513] = -'sd55016;
    data[ 1514] = -'sd57430;
    data[ 1515] = -'sd74328;
    data[ 1516] = -'sd28773;
    data[ 1517] = -'sd37570;
    data[ 1518] =  'sd64692;
    data[ 1519] = -'sd38679;
    data[ 1520] =  'sd56929;
    data[ 1521] =  'sd70821;
    data[ 1522] =  'sd4224;
    data[ 1523] =  'sd29568;
    data[ 1524] =  'sd43135;
    data[ 1525] = -'sd25737;
    data[ 1526] = -'sd16318;
    data[ 1527] =  'sd49615;
    data[ 1528] =  'sd19623;
    data[ 1529] = -'sd26480;
    data[ 1530] = -'sd21519;
    data[ 1531] =  'sd13208;
    data[ 1532] = -'sd71385;
    data[ 1533] = -'sd8172;
    data[ 1534] = -'sd57204;
    data[ 1535] = -'sd72746;
    data[ 1536] = -'sd17699;
    data[ 1537] =  'sd39948;
    data[ 1538] = -'sd48046;
    data[ 1539] = -'sd8640;
    data[ 1540] = -'sd60480;
    data[ 1541] =  'sd68163;
    data[ 1542] = -'sd14382;
    data[ 1543] =  'sd63167;
    data[ 1544] = -'sd49354;
    data[ 1545] = -'sd17796;
    data[ 1546] =  'sd39269;
    data[ 1547] = -'sd52799;
    data[ 1548] = -'sd41911;
    data[ 1549] =  'sd34305;
    data[ 1550] =  'sd76294;
    data[ 1551] =  'sd42535;
    data[ 1552] = -'sd29937;
    data[ 1553] = -'sd45718;
    data[ 1554] =  'sd7656;
    data[ 1555] =  'sd53592;
    data[ 1556] =  'sd47462;
    data[ 1557] =  'sd4552;
    data[ 1558] =  'sd31864;
    data[ 1559] =  'sd59207;
    data[ 1560] = -'sd77074;
    data[ 1561] = -'sd47995;
    data[ 1562] = -'sd8283;
    data[ 1563] = -'sd57981;
    data[ 1564] = -'sd78185;
    data[ 1565] = -'sd55772;
    data[ 1566] = -'sd62722;
    data[ 1567] =  'sd52469;
    data[ 1568] =  'sd39601;
    data[ 1569] = -'sd50475;
    data[ 1570] = -'sd25643;
    data[ 1571] = -'sd15660;
    data[ 1572] =  'sd54221;
    data[ 1573] =  'sd51865;
    data[ 1574] =  'sd35373;
    data[ 1575] = -'sd80071;
    data[ 1576] = -'sd68974;
    data[ 1577] =  'sd8705;
    data[ 1578] =  'sd60935;
    data[ 1579] = -'sd64978;
    data[ 1580] =  'sd36677;
    data[ 1581] = -'sd70943;
    data[ 1582] = -'sd5078;
    data[ 1583] = -'sd35546;
    data[ 1584] =  'sd78860;
    data[ 1585] =  'sd60497;
    data[ 1586] = -'sd68044;
    data[ 1587] =  'sd15215;
    data[ 1588] = -'sd57336;
    data[ 1589] = -'sd73670;
    data[ 1590] = -'sd24167;
    data[ 1591] = -'sd5328;
    data[ 1592] = -'sd37296;
    data[ 1593] =  'sd66610;
    data[ 1594] = -'sd25253;
    data[ 1595] = -'sd12930;
    data[ 1596] =  'sd73331;
    data[ 1597] =  'sd21794;
    data[ 1598] = -'sd11283;
    data[ 1599] = -'sd78981;
    data[ 1600] = -'sd61344;
    data[ 1601] =  'sd62115;
    data[ 1602] = -'sd56718;
    data[ 1603] = -'sd69344;
    data[ 1604] =  'sd6115;
    data[ 1605] =  'sd42805;
    data[ 1606] = -'sd28047;
    data[ 1607] = -'sd32488;
    data[ 1608] = -'sd63575;
    data[ 1609] =  'sd46498;
    data[ 1610] = -'sd2196;
    data[ 1611] = -'sd15372;
    data[ 1612] =  'sd56237;
    data[ 1613] =  'sd65977;
    data[ 1614] = -'sd29684;
    data[ 1615] = -'sd43947;
    data[ 1616] =  'sd20053;
    data[ 1617] = -'sd23470;
    data[ 1618] = -'sd449;
    data[ 1619] = -'sd3143;
    data[ 1620] = -'sd22001;
    data[ 1621] =  'sd9834;
    data[ 1622] =  'sd68838;
    data[ 1623] = -'sd9657;
    data[ 1624] = -'sd67599;
    data[ 1625] =  'sd18330;
    data[ 1626] = -'sd35531;
    data[ 1627] =  'sd78965;
    data[ 1628] =  'sd61232;
    data[ 1629] = -'sd62899;
    data[ 1630] =  'sd51230;
    data[ 1631] =  'sd30928;
    data[ 1632] =  'sd52655;
    data[ 1633] =  'sd40903;
    data[ 1634] = -'sd41361;
    data[ 1635] =  'sd38155;
    data[ 1636] = -'sd60597;
    data[ 1637] =  'sd67344;
    data[ 1638] = -'sd20115;
    data[ 1639] =  'sd23036;
    data[ 1640] = -'sd2589;
    data[ 1641] = -'sd18123;
    data[ 1642] =  'sd36980;
    data[ 1643] = -'sd68822;
    data[ 1644] =  'sd9769;
    data[ 1645] =  'sd68383;
    data[ 1646] = -'sd12842;
    data[ 1647] =  'sd73947;
    data[ 1648] =  'sd26106;
    data[ 1649] =  'sd18901;
    data[ 1650] = -'sd31534;
    data[ 1651] = -'sd56897;
    data[ 1652] = -'sd70597;
    data[ 1653] = -'sd2656;
    data[ 1654] = -'sd18592;
    data[ 1655] =  'sd33697;
    data[ 1656] =  'sd72038;
    data[ 1657] =  'sd12743;
    data[ 1658] = -'sd74640;
    data[ 1659] = -'sd30957;
    data[ 1660] = -'sd52858;
    data[ 1661] = -'sd42324;
    data[ 1662] =  'sd31414;
    data[ 1663] =  'sd56057;
    data[ 1664] =  'sd64717;
    data[ 1665] = -'sd38504;
    data[ 1666] =  'sd58154;
    data[ 1667] =  'sd79396;
    data[ 1668] =  'sd64249;
    data[ 1669] = -'sd41780;
    data[ 1670] =  'sd35222;
    data[ 1671] = -'sd81128;
    data[ 1672] = -'sd76373;
    data[ 1673] = -'sd43088;
    data[ 1674] =  'sd26066;
    data[ 1675] =  'sd18621;
    data[ 1676] = -'sd33494;
    data[ 1677] = -'sd70617;
    data[ 1678] = -'sd2796;
    data[ 1679] = -'sd19572;
    data[ 1680] =  'sd26837;
    data[ 1681] =  'sd24018;
    data[ 1682] =  'sd4285;
    data[ 1683] =  'sd29995;
    data[ 1684] =  'sd46124;
    data[ 1685] = -'sd4814;
    data[ 1686] = -'sd33698;
    data[ 1687] = -'sd72045;
    data[ 1688] = -'sd12792;
    data[ 1689] =  'sd74297;
    data[ 1690] =  'sd28556;
    data[ 1691] =  'sd36051;
    data[ 1692] = -'sd75325;
    data[ 1693] = -'sd35752;
    data[ 1694] =  'sd77418;
    data[ 1695] =  'sd50403;
    data[ 1696] =  'sd25139;
    data[ 1697] =  'sd12132;
    data[ 1698] = -'sd78917;
    data[ 1699] = -'sd60896;
    data[ 1700] =  'sd65251;
    data[ 1701] = -'sd34766;
    data[ 1702] = -'sd79521;
    data[ 1703] = -'sd65124;
    data[ 1704] =  'sd35655;
    data[ 1705] = -'sd78097;
    data[ 1706] = -'sd55156;
    data[ 1707] = -'sd58410;
    data[ 1708] = -'sd81188;
    data[ 1709] = -'sd76793;
    data[ 1710] = -'sd46028;
    data[ 1711] =  'sd5486;
    data[ 1712] =  'sd38402;
    data[ 1713] = -'sd58868;
    data[ 1714] =  'sd79447;
    data[ 1715] =  'sd64606;
    data[ 1716] = -'sd39281;
    data[ 1717] =  'sd52715;
    data[ 1718] =  'sd41323;
    data[ 1719] = -'sd38421;
    data[ 1720] =  'sd58735;
    data[ 1721] = -'sd80378;
    data[ 1722] = -'sd71123;
    data[ 1723] = -'sd6338;
    data[ 1724] = -'sd44366;
    data[ 1725] =  'sd17120;
    data[ 1726] = -'sd44001;
    data[ 1727] =  'sd19675;
    data[ 1728] = -'sd26116;
    data[ 1729] = -'sd18971;
    data[ 1730] =  'sd31044;
    data[ 1731] =  'sd53467;
    data[ 1732] =  'sd46587;
    data[ 1733] = -'sd1573;
    data[ 1734] = -'sd11011;
    data[ 1735] = -'sd77077;
    data[ 1736] = -'sd48016;
    data[ 1737] = -'sd8430;
    data[ 1738] = -'sd59010;
    data[ 1739] =  'sd78453;
    data[ 1740] =  'sd57648;
    data[ 1741] =  'sd75854;
    data[ 1742] =  'sd39455;
    data[ 1743] = -'sd51497;
    data[ 1744] = -'sd32797;
    data[ 1745] = -'sd65738;
    data[ 1746] =  'sd31357;
    data[ 1747] =  'sd55658;
    data[ 1748] =  'sd61924;
    data[ 1749] = -'sd58055;
    data[ 1750] = -'sd78703;
    data[ 1751] = -'sd59398;
    data[ 1752] =  'sd75737;
    data[ 1753] =  'sd38636;
    data[ 1754] = -'sd57230;
    data[ 1755] = -'sd72928;
    data[ 1756] = -'sd18973;
    data[ 1757] =  'sd31030;
    data[ 1758] =  'sd53369;
    data[ 1759] =  'sd45901;
    data[ 1760] = -'sd6375;
    data[ 1761] = -'sd44625;
    data[ 1762] =  'sd15307;
    data[ 1763] = -'sd56692;
    data[ 1764] = -'sd69162;
    data[ 1765] =  'sd7389;
    data[ 1766] =  'sd51723;
    data[ 1767] =  'sd34379;
    data[ 1768] =  'sd76812;
    data[ 1769] =  'sd46161;
    data[ 1770] = -'sd4555;
    data[ 1771] = -'sd31885;
    data[ 1772] = -'sd59354;
    data[ 1773] =  'sd76045;
    data[ 1774] =  'sd40792;
    data[ 1775] = -'sd42138;
    data[ 1776] =  'sd32716;
    data[ 1777] =  'sd65171;
    data[ 1778] = -'sd35326;
    data[ 1779] =  'sd80400;
    data[ 1780] =  'sd71277;
    data[ 1781] =  'sd7416;
    data[ 1782] =  'sd51912;
    data[ 1783] =  'sd35702;
    data[ 1784] = -'sd77768;
    data[ 1785] = -'sd52853;
    data[ 1786] = -'sd42289;
    data[ 1787] =  'sd31659;
    data[ 1788] =  'sd57772;
    data[ 1789] =  'sd76722;
    data[ 1790] =  'sd45531;
    data[ 1791] = -'sd8965;
    data[ 1792] = -'sd62755;
    data[ 1793] =  'sd52238;
    data[ 1794] =  'sd37984;
    data[ 1795] = -'sd61794;
    data[ 1796] =  'sd58965;
    data[ 1797] = -'sd78768;
    data[ 1798] = -'sd59853;
    data[ 1799] =  'sd72552;
    data[ 1800] =  'sd16341;
    data[ 1801] = -'sd49454;
    data[ 1802] = -'sd18496;
    data[ 1803] =  'sd34369;
    data[ 1804] =  'sd76742;
    data[ 1805] =  'sd45671;
    data[ 1806] = -'sd7985;
    data[ 1807] = -'sd55895;
    data[ 1808] = -'sd63583;
    data[ 1809] =  'sd46442;
    data[ 1810] = -'sd2588;
    data[ 1811] = -'sd18116;
    data[ 1812] =  'sd37029;
    data[ 1813] = -'sd68479;
    data[ 1814] =  'sd12170;
    data[ 1815] = -'sd78651;
    data[ 1816] = -'sd59034;
    data[ 1817] =  'sd78285;
    data[ 1818] =  'sd56472;
    data[ 1819] =  'sd67622;
    data[ 1820] = -'sd18169;
    data[ 1821] =  'sd36658;
    data[ 1822] = -'sd71076;
    data[ 1823] = -'sd6009;
    data[ 1824] = -'sd42063;
    data[ 1825] =  'sd33241;
    data[ 1826] =  'sd68846;
    data[ 1827] = -'sd9601;
    data[ 1828] = -'sd67207;
    data[ 1829] =  'sd21074;
    data[ 1830] = -'sd16323;
    data[ 1831] =  'sd49580;
    data[ 1832] =  'sd19378;
    data[ 1833] = -'sd28195;
    data[ 1834] = -'sd33524;
    data[ 1835] = -'sd70827;
    data[ 1836] = -'sd4266;
    data[ 1837] = -'sd29862;
    data[ 1838] = -'sd45193;
    data[ 1839] =  'sd11331;
    data[ 1840] =  'sd79317;
    data[ 1841] =  'sd63696;
    data[ 1842] = -'sd45651;
    data[ 1843] =  'sd8125;
    data[ 1844] =  'sd56875;
    data[ 1845] =  'sd70443;
    data[ 1846] =  'sd1578;
    data[ 1847] =  'sd11046;
    data[ 1848] =  'sd77322;
    data[ 1849] =  'sd49731;
    data[ 1850] =  'sd20435;
    data[ 1851] = -'sd20796;
    data[ 1852] =  'sd18269;
    data[ 1853] = -'sd35958;
    data[ 1854] =  'sd75976;
    data[ 1855] =  'sd40309;
    data[ 1856] = -'sd45519;
    data[ 1857] =  'sd9049;
    data[ 1858] =  'sd63343;
    data[ 1859] = -'sd48122;
    data[ 1860] = -'sd9172;
    data[ 1861] = -'sd64204;
    data[ 1862] =  'sd42095;
    data[ 1863] = -'sd33017;
    data[ 1864] = -'sd67278;
    data[ 1865] =  'sd20577;
    data[ 1866] = -'sd19802;
    data[ 1867] =  'sd25227;
    data[ 1868] =  'sd12748;
    data[ 1869] = -'sd74605;
    data[ 1870] = -'sd30712;
    data[ 1871] = -'sd51143;
    data[ 1872] = -'sd30319;
    data[ 1873] = -'sd48392;
    data[ 1874] = -'sd11062;
    data[ 1875] = -'sd77434;
    data[ 1876] = -'sd50515;
    data[ 1877] = -'sd25923;
    data[ 1878] = -'sd17620;
    data[ 1879] =  'sd40501;
    data[ 1880] = -'sd44175;
    data[ 1881] =  'sd18457;
    data[ 1882] = -'sd34642;
    data[ 1883] = -'sd78653;
    data[ 1884] = -'sd59048;
    data[ 1885] =  'sd78187;
    data[ 1886] =  'sd55786;
    data[ 1887] =  'sd62820;
    data[ 1888] = -'sd51783;
    data[ 1889] = -'sd34799;
    data[ 1890] = -'sd79752;
    data[ 1891] = -'sd66741;
    data[ 1892] =  'sd24336;
    data[ 1893] =  'sd6511;
    data[ 1894] =  'sd45577;
    data[ 1895] = -'sd8643;
    data[ 1896] = -'sd60501;
    data[ 1897] =  'sd68016;
    data[ 1898] = -'sd15411;
    data[ 1899] =  'sd55964;
    data[ 1900] =  'sd64066;
    data[ 1901] = -'sd43061;
    data[ 1902] =  'sd26255;
    data[ 1903] =  'sd19944;
    data[ 1904] = -'sd24233;
    data[ 1905] = -'sd5790;
    data[ 1906] = -'sd40530;
    data[ 1907] =  'sd43972;
    data[ 1908] = -'sd19878;
    data[ 1909] =  'sd24695;
    data[ 1910] =  'sd9024;
    data[ 1911] =  'sd63168;
    data[ 1912] = -'sd49347;
    data[ 1913] = -'sd17747;
    data[ 1914] =  'sd39612;
    data[ 1915] = -'sd50398;
    data[ 1916] = -'sd25104;
    data[ 1917] = -'sd11887;
    data[ 1918] =  'sd80632;
    data[ 1919] =  'sd72901;
    data[ 1920] =  'sd18784;
    data[ 1921] = -'sd32353;
    data[ 1922] = -'sd62630;
    data[ 1923] =  'sd53113;
    data[ 1924] =  'sd44109;
    data[ 1925] = -'sd18919;
    data[ 1926] =  'sd31408;
    data[ 1927] =  'sd56015;
    data[ 1928] =  'sd64423;
    data[ 1929] = -'sd40562;
    data[ 1930] =  'sd43748;
    data[ 1931] = -'sd21446;
    data[ 1932] =  'sd13719;
    data[ 1933] = -'sd67808;
    data[ 1934] =  'sd16867;
    data[ 1935] = -'sd45772;
    data[ 1936] =  'sd7278;
    data[ 1937] =  'sd50946;
    data[ 1938] =  'sd28940;
    data[ 1939] =  'sd38739;
    data[ 1940] = -'sd56509;
    data[ 1941] = -'sd67881;
    data[ 1942] =  'sd16356;
    data[ 1943] = -'sd49349;
    data[ 1944] = -'sd17761;
    data[ 1945] =  'sd39514;
    data[ 1946] = -'sd51084;
    data[ 1947] = -'sd29906;
    data[ 1948] = -'sd45501;
    data[ 1949] =  'sd9175;
    data[ 1950] =  'sd64225;
    data[ 1951] = -'sd41948;
    data[ 1952] =  'sd34046;
    data[ 1953] =  'sd74481;
    data[ 1954] =  'sd29844;
    data[ 1955] =  'sd45067;
    data[ 1956] = -'sd12213;
    data[ 1957] =  'sd78350;
    data[ 1958] =  'sd56927;
    data[ 1959] =  'sd70807;
    data[ 1960] =  'sd4126;
    data[ 1961] =  'sd28882;
    data[ 1962] =  'sd38333;
    data[ 1963] = -'sd59351;
    data[ 1964] =  'sd76066;
    data[ 1965] =  'sd40939;
    data[ 1966] = -'sd41109;
    data[ 1967] =  'sd39919;
    data[ 1968] = -'sd48249;
    data[ 1969] = -'sd10061;
    data[ 1970] = -'sd70427;
    data[ 1971] = -'sd1466;
    data[ 1972] = -'sd10262;
    data[ 1973] = -'sd71834;
    data[ 1974] = -'sd11315;
    data[ 1975] = -'sd79205;
    data[ 1976] = -'sd62912;
    data[ 1977] =  'sd51139;
    data[ 1978] =  'sd30291;
    data[ 1979] =  'sd48196;
    data[ 1980] =  'sd9690;
    data[ 1981] =  'sd67830;
    data[ 1982] = -'sd16713;
    data[ 1983] =  'sd46850;
    data[ 1984] =  'sd268;
    data[ 1985] =  'sd1876;
    data[ 1986] =  'sd13132;
    data[ 1987] = -'sd71917;
    data[ 1988] = -'sd11896;
    data[ 1989] =  'sd80569;
    data[ 1990] =  'sd72460;
    data[ 1991] =  'sd15697;
    data[ 1992] = -'sd53962;
    data[ 1993] = -'sd50052;
    data[ 1994] = -'sd22682;
    data[ 1995] =  'sd5067;
    data[ 1996] =  'sd35469;
    data[ 1997] = -'sd79399;
    data[ 1998] = -'sd64270;
    data[ 1999] =  'sd41633;
    data[ 2000] = -'sd36251;
    data[ 2001] =  'sd73925;
    data[ 2002] =  'sd25952;
    data[ 2003] =  'sd17823;
    data[ 2004] = -'sd39080;
    data[ 2005] =  'sd54122;
    data[ 2006] =  'sd51172;
    data[ 2007] =  'sd30522;
    data[ 2008] =  'sd49813;
    data[ 2009] =  'sd21009;
    data[ 2010] = -'sd16778;
    data[ 2011] =  'sd46395;
    data[ 2012] = -'sd2917;
    data[ 2013] = -'sd20419;
    data[ 2014] =  'sd20908;
    data[ 2015] = -'sd17485;
    data[ 2016] =  'sd41446;
    data[ 2017] = -'sd37560;
    data[ 2018] =  'sd64762;
    data[ 2019] = -'sd38189;
    data[ 2020] =  'sd60359;
    data[ 2021] = -'sd69010;
    data[ 2022] =  'sd8453;
    data[ 2023] =  'sd59171;
    data[ 2024] = -'sd77326;
    data[ 2025] = -'sd49759;
    data[ 2026] = -'sd20631;
    data[ 2027] =  'sd19424;
    data[ 2028] = -'sd27873;
    data[ 2029] = -'sd31270;
    data[ 2030] = -'sd55049;
    data[ 2031] = -'sd57661;
    data[ 2032] = -'sd75945;
    data[ 2033] = -'sd40092;
    data[ 2034] =  'sd47038;
    data[ 2035] =  'sd1584;
    data[ 2036] =  'sd11088;
    data[ 2037] =  'sd77616;
    data[ 2038] =  'sd51789;
    data[ 2039] =  'sd34841;
    data[ 2040] =  'sd80046;
    data[ 2041] =  'sd68799;
    data[ 2042] = -'sd9930;
    data[ 2043] = -'sd69510;
    data[ 2044] =  'sd4953;
    data[ 2045] =  'sd34671;
    data[ 2046] =  'sd78856;
    data[ 2047] =  'sd60469;
    data[ 2048] = -'sd68240;
    data[ 2049] =  'sd13843;
    data[ 2050] = -'sd66940;
    data[ 2051] =  'sd22943;
    data[ 2052] = -'sd3240;
    data[ 2053] = -'sd22680;
    data[ 2054] =  'sd5081;
    data[ 2055] =  'sd35567;
    data[ 2056] = -'sd78713;
    data[ 2057] = -'sd59468;
    data[ 2058] =  'sd75247;
    data[ 2059] =  'sd35206;
    data[ 2060] = -'sd81240;
    data[ 2061] = -'sd77157;
    data[ 2062] = -'sd48576;
    data[ 2063] = -'sd12350;
    data[ 2064] =  'sd77391;
    data[ 2065] =  'sd50214;
    data[ 2066] =  'sd23816;
    data[ 2067] =  'sd2871;
    data[ 2068] =  'sd20097;
    data[ 2069] = -'sd23162;
    data[ 2070] =  'sd1707;
    data[ 2071] =  'sd11949;
    data[ 2072] = -'sd80198;
    data[ 2073] = -'sd69863;
    data[ 2074] =  'sd2482;
    data[ 2075] =  'sd17374;
    data[ 2076] = -'sd42223;
    data[ 2077] =  'sd32121;
    data[ 2078] =  'sd61006;
    data[ 2079] = -'sd64481;
    data[ 2080] =  'sd40156;
    data[ 2081] = -'sd46590;
    data[ 2082] =  'sd1552;
    data[ 2083] =  'sd10864;
    data[ 2084] =  'sd76048;
    data[ 2085] =  'sd40813;
    data[ 2086] = -'sd41991;
    data[ 2087] =  'sd33745;
    data[ 2088] =  'sd72374;
    data[ 2089] =  'sd15095;
    data[ 2090] = -'sd58176;
    data[ 2091] = -'sd79550;
    data[ 2092] = -'sd65327;
    data[ 2093] =  'sd34234;
    data[ 2094] =  'sd75797;
    data[ 2095] =  'sd39056;
    data[ 2096] = -'sd54290;
    data[ 2097] = -'sd52348;
    data[ 2098] = -'sd38754;
    data[ 2099] =  'sd56404;
    data[ 2100] =  'sd67146;
    data[ 2101] = -'sd21501;
    data[ 2102] =  'sd13334;
    data[ 2103] = -'sd70503;
    data[ 2104] = -'sd1998;
    data[ 2105] = -'sd13986;
    data[ 2106] =  'sd65939;
    data[ 2107] = -'sd29950;
    data[ 2108] = -'sd45809;
    data[ 2109] =  'sd7019;
    data[ 2110] =  'sd49133;
    data[ 2111] =  'sd16249;
    data[ 2112] = -'sd50098;
    data[ 2113] = -'sd23004;
    data[ 2114] =  'sd2813;
    data[ 2115] =  'sd19691;
    data[ 2116] = -'sd26004;
    data[ 2117] = -'sd18187;
    data[ 2118] =  'sd36532;
    data[ 2119] = -'sd71958;
    data[ 2120] = -'sd12183;
    data[ 2121] =  'sd78560;
    data[ 2122] =  'sd58397;
    data[ 2123] =  'sd81097;
    data[ 2124] =  'sd76156;
    data[ 2125] =  'sd41569;
    data[ 2126] = -'sd36699;
    data[ 2127] =  'sd70789;
    data[ 2128] =  'sd4000;
    data[ 2129] =  'sd28000;
    data[ 2130] =  'sd32159;
    data[ 2131] =  'sd61272;
    data[ 2132] = -'sd62619;
    data[ 2133] =  'sd53190;
    data[ 2134] =  'sd44648;
    data[ 2135] = -'sd15146;
    data[ 2136] =  'sd57819;
    data[ 2137] =  'sd77051;
    data[ 2138] =  'sd47834;
    data[ 2139] =  'sd7156;
    data[ 2140] =  'sd50092;
    data[ 2141] =  'sd22962;
    data[ 2142] = -'sd3107;
    data[ 2143] = -'sd21749;
    data[ 2144] =  'sd11598;
    data[ 2145] =  'sd81186;
    data[ 2146] =  'sd76779;
    data[ 2147] =  'sd45930;
    data[ 2148] = -'sd6172;
    data[ 2149] = -'sd43204;
    data[ 2150] =  'sd25254;
    data[ 2151] =  'sd12937;
    data[ 2152] = -'sd73282;
    data[ 2153] = -'sd21451;
    data[ 2154] =  'sd13684;
    data[ 2155] = -'sd68053;
    data[ 2156] =  'sd15152;
    data[ 2157] = -'sd57777;
    data[ 2158] = -'sd76757;
    data[ 2159] = -'sd45776;
    data[ 2160] =  'sd7250;
    data[ 2161] =  'sd50750;
    data[ 2162] =  'sd27568;
    data[ 2163] =  'sd29135;
    data[ 2164] =  'sd40104;
    data[ 2165] = -'sd46954;
    data[ 2166] = -'sd996;
    data[ 2167] = -'sd6972;
    data[ 2168] = -'sd48804;
    data[ 2169] = -'sd13946;
    data[ 2170] =  'sd66219;
    data[ 2171] = -'sd27990;
    data[ 2172] = -'sd32089;
    data[ 2173] = -'sd60782;
    data[ 2174] =  'sd66049;
    data[ 2175] = -'sd29180;
    data[ 2176] = -'sd40419;
    data[ 2177] =  'sd44749;
    data[ 2178] = -'sd14439;
    data[ 2179] =  'sd62768;
    data[ 2180] = -'sd52147;
    data[ 2181] = -'sd37347;
    data[ 2182] =  'sd66253;
    data[ 2183] = -'sd27752;
    data[ 2184] = -'sd30423;
    data[ 2185] = -'sd49120;
    data[ 2186] = -'sd16158;
    data[ 2187] =  'sd50735;
    data[ 2188] =  'sd27463;
    data[ 2189] =  'sd28400;
    data[ 2190] =  'sd34959;
    data[ 2191] =  'sd80872;
    data[ 2192] =  'sd74581;
    data[ 2193] =  'sd30544;
    data[ 2194] =  'sd49967;
    data[ 2195] =  'sd22087;
    data[ 2196] = -'sd9232;
    data[ 2197] = -'sd64624;
    data[ 2198] =  'sd39155;
    data[ 2199] = -'sd53597;
    data[ 2200] = -'sd47497;
    data[ 2201] = -'sd4797;
    data[ 2202] = -'sd33579;
    data[ 2203] = -'sd71212;
    data[ 2204] = -'sd6961;
    data[ 2205] = -'sd48727;
    data[ 2206] = -'sd13407;
    data[ 2207] =  'sd69992;
    data[ 2208] = -'sd1579;
    data[ 2209] = -'sd11053;
    data[ 2210] = -'sd77371;
    data[ 2211] = -'sd50074;
    data[ 2212] = -'sd22836;
    data[ 2213] =  'sd3989;
    data[ 2214] =  'sd27923;
    data[ 2215] =  'sd31620;
    data[ 2216] =  'sd57499;
    data[ 2217] =  'sd74811;
    data[ 2218] =  'sd32154;
    data[ 2219] =  'sd61237;
    data[ 2220] = -'sd62864;
    data[ 2221] =  'sd51475;
    data[ 2222] =  'sd32643;
    data[ 2223] =  'sd64660;
    data[ 2224] = -'sd38903;
    data[ 2225] =  'sd55361;
    data[ 2226] =  'sd59845;
    data[ 2227] = -'sd72608;
    data[ 2228] = -'sd16733;
    data[ 2229] =  'sd46710;
    data[ 2230] = -'sd712;
    data[ 2231] = -'sd4984;
    data[ 2232] = -'sd34888;
    data[ 2233] = -'sd80375;
    data[ 2234] = -'sd71102;
    data[ 2235] = -'sd6191;
    data[ 2236] = -'sd43337;
    data[ 2237] =  'sd24323;
    data[ 2238] =  'sd6420;
    data[ 2239] =  'sd44940;
    data[ 2240] = -'sd13102;
    data[ 2241] =  'sd72127;
    data[ 2242] =  'sd13366;
    data[ 2243] = -'sd70279;
    data[ 2244] = -'sd430;
    data[ 2245] = -'sd3010;
    data[ 2246] = -'sd21070;
    data[ 2247] =  'sd16351;
    data[ 2248] = -'sd49384;
    data[ 2249] = -'sd18006;
    data[ 2250] =  'sd37799;
    data[ 2251] = -'sd63089;
    data[ 2252] =  'sd49900;
    data[ 2253] =  'sd21618;
    data[ 2254] = -'sd12515;
    data[ 2255] =  'sd76236;
    data[ 2256] =  'sd42129;
    data[ 2257] = -'sd32779;
    data[ 2258] = -'sd65612;
    data[ 2259] =  'sd32239;
    data[ 2260] =  'sd61832;
    data[ 2261] = -'sd58699;
    data[ 2262] =  'sd80630;
    data[ 2263] =  'sd72887;
    data[ 2264] =  'sd18686;
    data[ 2265] = -'sd33039;
    data[ 2266] = -'sd67432;
    data[ 2267] =  'sd19499;
    data[ 2268] = -'sd27348;
    data[ 2269] = -'sd27595;
    data[ 2270] = -'sd29324;
    data[ 2271] = -'sd41427;
    data[ 2272] =  'sd37693;
    data[ 2273] = -'sd63831;
    data[ 2274] =  'sd44706;
    data[ 2275] = -'sd14740;
    data[ 2276] =  'sd60661;
    data[ 2277] = -'sd66896;
    data[ 2278] =  'sd23251;
    data[ 2279] = -'sd1084;
    data[ 2280] = -'sd7588;
    data[ 2281] = -'sd53116;
    data[ 2282] = -'sd44130;
    data[ 2283] =  'sd18772;
    data[ 2284] = -'sd32437;
    data[ 2285] = -'sd63218;
    data[ 2286] =  'sd48997;
    data[ 2287] =  'sd15297;
    data[ 2288] = -'sd56762;
    data[ 2289] = -'sd69652;
    data[ 2290] =  'sd3959;
    data[ 2291] =  'sd27713;
    data[ 2292] =  'sd30150;
    data[ 2293] =  'sd47209;
    data[ 2294] =  'sd2781;
    data[ 2295] =  'sd19467;
    data[ 2296] = -'sd27572;
    data[ 2297] = -'sd29163;
    data[ 2298] = -'sd40300;
    data[ 2299] =  'sd45582;
    data[ 2300] = -'sd8608;
    data[ 2301] = -'sd60256;
    data[ 2302] =  'sd69731;
    data[ 2303] = -'sd3406;
    data[ 2304] = -'sd23842;
    data[ 2305] = -'sd3053;
    data[ 2306] = -'sd21371;
    data[ 2307] =  'sd14244;
    data[ 2308] = -'sd64133;
    data[ 2309] =  'sd42592;
    data[ 2310] = -'sd29538;
    data[ 2311] = -'sd42925;
    data[ 2312] =  'sd27207;
    data[ 2313] =  'sd26608;
    data[ 2314] =  'sd22415;
    data[ 2315] = -'sd6936;
    data[ 2316] = -'sd48552;
    data[ 2317] = -'sd12182;
    data[ 2318] =  'sd78567;
    data[ 2319] =  'sd58446;
    data[ 2320] =  'sd81440;
    data[ 2321] =  'sd78557;
    data[ 2322] =  'sd58376;
    data[ 2323] =  'sd80950;
    data[ 2324] =  'sd75127;
    data[ 2325] =  'sd34366;
    data[ 2326] =  'sd76721;
    data[ 2327] =  'sd45524;
    data[ 2328] = -'sd9014;
    data[ 2329] = -'sd63098;
    data[ 2330] =  'sd49837;
    data[ 2331] =  'sd21177;
    data[ 2332] = -'sd15602;
    data[ 2333] =  'sd54627;
    data[ 2334] =  'sd54707;
    data[ 2335] =  'sd55267;
    data[ 2336] =  'sd59187;
    data[ 2337] = -'sd77214;
    data[ 2338] = -'sd48975;
    data[ 2339] = -'sd15143;
    data[ 2340] =  'sd57840;
    data[ 2341] =  'sd77198;
    data[ 2342] =  'sd48863;
    data[ 2343] =  'sd14359;
    data[ 2344] = -'sd63328;
    data[ 2345] =  'sd48227;
    data[ 2346] =  'sd9907;
    data[ 2347] =  'sd69349;
    data[ 2348] = -'sd6080;
    data[ 2349] = -'sd42560;
    data[ 2350] =  'sd29762;
    data[ 2351] =  'sd44493;
    data[ 2352] = -'sd16231;
    data[ 2353] =  'sd50224;
    data[ 2354] =  'sd23886;
    data[ 2355] =  'sd3361;
    data[ 2356] =  'sd23527;
    data[ 2357] =  'sd848;
    data[ 2358] =  'sd5936;
    data[ 2359] =  'sd41552;
    data[ 2360] = -'sd36818;
    data[ 2361] =  'sd69956;
    data[ 2362] = -'sd1831;
    data[ 2363] = -'sd12817;
    data[ 2364] =  'sd74122;
    data[ 2365] =  'sd27331;
    data[ 2366] =  'sd27476;
    data[ 2367] =  'sd28491;
    data[ 2368] =  'sd35596;
    data[ 2369] = -'sd78510;
    data[ 2370] = -'sd58047;
    data[ 2371] = -'sd78647;
    data[ 2372] = -'sd59006;
    data[ 2373] =  'sd78481;
    data[ 2374] =  'sd57844;
    data[ 2375] =  'sd77226;
    data[ 2376] =  'sd49059;
    data[ 2377] =  'sd15731;
    data[ 2378] = -'sd53724;
    data[ 2379] = -'sd48386;
    data[ 2380] = -'sd11020;
    data[ 2381] = -'sd77140;
    data[ 2382] = -'sd48457;
    data[ 2383] = -'sd11517;
    data[ 2384] = -'sd80619;
    data[ 2385] = -'sd72810;
    data[ 2386] = -'sd18147;
    data[ 2387] =  'sd36812;
    data[ 2388] = -'sd69998;
    data[ 2389] =  'sd1537;
    data[ 2390] =  'sd10759;
    data[ 2391] =  'sd75313;
    data[ 2392] =  'sd35668;
    data[ 2393] = -'sd78006;
    data[ 2394] = -'sd54519;
    data[ 2395] = -'sd53951;
    data[ 2396] = -'sd49975;
    data[ 2397] = -'sd22143;
    data[ 2398] =  'sd8840;
    data[ 2399] =  'sd61880;
    data[ 2400] = -'sd58363;
    data[ 2401] = -'sd80859;
    data[ 2402] = -'sd74490;
    data[ 2403] = -'sd29907;
    data[ 2404] = -'sd45508;
    data[ 2405] =  'sd9126;
    data[ 2406] =  'sd63882;
    data[ 2407] = -'sd44349;
    data[ 2408] =  'sd17239;
    data[ 2409] = -'sd43168;
    data[ 2410] =  'sd25506;
    data[ 2411] =  'sd14701;
    data[ 2412] = -'sd60934;
    data[ 2413] =  'sd64985;
    data[ 2414] = -'sd36628;
    data[ 2415] =  'sd71286;
    data[ 2416] =  'sd7479;
    data[ 2417] =  'sd52353;
    data[ 2418] =  'sd38789;
    data[ 2419] = -'sd56159;
    data[ 2420] = -'sd65431;
    data[ 2421] =  'sd33506;
    data[ 2422] =  'sd70701;
    data[ 2423] =  'sd3384;
    data[ 2424] =  'sd23688;
    data[ 2425] =  'sd1975;
    data[ 2426] =  'sd13825;
    data[ 2427] = -'sd67066;
    data[ 2428] =  'sd22061;
    data[ 2429] = -'sd9414;
    data[ 2430] = -'sd65898;
    data[ 2431] =  'sd30237;
    data[ 2432] =  'sd47818;
    data[ 2433] =  'sd7044;
    data[ 2434] =  'sd49308;
    data[ 2435] =  'sd17474;
    data[ 2436] = -'sd41523;
    data[ 2437] =  'sd37021;
    data[ 2438] = -'sd68535;
    data[ 2439] =  'sd11778;
    data[ 2440] = -'sd81395;
    data[ 2441] = -'sd78242;
    data[ 2442] = -'sd56171;
    data[ 2443] = -'sd65515;
    data[ 2444] =  'sd32918;
    data[ 2445] =  'sd66585;
    data[ 2446] = -'sd25428;
    data[ 2447] = -'sd14155;
    data[ 2448] =  'sd64756;
    data[ 2449] = -'sd38231;
    data[ 2450] =  'sd60065;
    data[ 2451] = -'sd71068;
    data[ 2452] = -'sd5953;
    data[ 2453] = -'sd41671;
    data[ 2454] =  'sd35985;
    data[ 2455] = -'sd75787;
    data[ 2456] = -'sd38986;
    data[ 2457] =  'sd54780;
    data[ 2458] =  'sd55778;
    data[ 2459] =  'sd62764;
    data[ 2460] = -'sd52175;
    data[ 2461] = -'sd37543;
    data[ 2462] =  'sd64881;
    data[ 2463] = -'sd37356;
    data[ 2464] =  'sd66190;
    data[ 2465] = -'sd28193;
    data[ 2466] = -'sd33510;
    data[ 2467] = -'sd70729;
    data[ 2468] = -'sd3580;
    data[ 2469] = -'sd25060;
    data[ 2470] = -'sd11579;
    data[ 2471] = -'sd81053;
    data[ 2472] = -'sd75848;
    data[ 2473] = -'sd39413;
    data[ 2474] =  'sd51791;
    data[ 2475] =  'sd34855;
    data[ 2476] =  'sd80144;
    data[ 2477] =  'sd69485;
    data[ 2478] = -'sd5128;
    data[ 2479] = -'sd35896;
    data[ 2480] =  'sd76410;
    data[ 2481] =  'sd43347;
    data[ 2482] = -'sd24253;
    data[ 2483] = -'sd5930;
    data[ 2484] = -'sd41510;
    data[ 2485] =  'sd37112;
    data[ 2486] = -'sd67898;
    data[ 2487] =  'sd16237;
    data[ 2488] = -'sd50182;
    data[ 2489] = -'sd23592;
    data[ 2490] = -'sd1303;
    data[ 2491] = -'sd9121;
    data[ 2492] = -'sd63847;
    data[ 2493] =  'sd44594;
    data[ 2494] = -'sd15524;
    data[ 2495] =  'sd55173;
    data[ 2496] =  'sd58529;
    data[ 2497] = -'sd81820;
    data[ 2498] = -'sd81217;
    data[ 2499] = -'sd76996;
    data[ 2500] = -'sd47449;
    data[ 2501] = -'sd4461;
    data[ 2502] = -'sd31227;
    data[ 2503] = -'sd54748;
    data[ 2504] = -'sd55554;
    data[ 2505] = -'sd61196;
    data[ 2506] =  'sd63151;
    data[ 2507] = -'sd49466;
    data[ 2508] = -'sd18580;
    data[ 2509] =  'sd33781;
    data[ 2510] =  'sd72626;
    data[ 2511] =  'sd16859;
    data[ 2512] = -'sd45828;
    data[ 2513] =  'sd6886;
    data[ 2514] =  'sd48202;
    data[ 2515] =  'sd9732;
    data[ 2516] =  'sd68124;
    data[ 2517] = -'sd14655;
    data[ 2518] =  'sd61256;
    data[ 2519] = -'sd62731;
    data[ 2520] =  'sd52406;
    data[ 2521] =  'sd39160;
    data[ 2522] = -'sd53562;
    data[ 2523] = -'sd47252;
    data[ 2524] = -'sd3082;
    data[ 2525] = -'sd21574;
    data[ 2526] =  'sd12823;
    data[ 2527] = -'sd74080;
    data[ 2528] = -'sd27037;
    data[ 2529] = -'sd25418;
    data[ 2530] = -'sd14085;
    data[ 2531] =  'sd65246;
    data[ 2532] = -'sd34801;
    data[ 2533] = -'sd79766;
    data[ 2534] = -'sd66839;
    data[ 2535] =  'sd23650;
    data[ 2536] =  'sd1709;
    data[ 2537] =  'sd11963;
    data[ 2538] = -'sd80100;
    data[ 2539] = -'sd69177;
    data[ 2540] =  'sd7284;
    data[ 2541] =  'sd50988;
    data[ 2542] =  'sd29234;
    data[ 2543] =  'sd40797;
    data[ 2544] = -'sd42103;
    data[ 2545] =  'sd32961;
    data[ 2546] =  'sd66886;
    data[ 2547] = -'sd23321;
    data[ 2548] =  'sd594;
    data[ 2549] =  'sd4158;
    data[ 2550] =  'sd29106;
    data[ 2551] =  'sd39901;
    data[ 2552] = -'sd48375;
    data[ 2553] = -'sd10943;
    data[ 2554] = -'sd76601;
    data[ 2555] = -'sd44684;
    data[ 2556] =  'sd14894;
    data[ 2557] = -'sd59583;
    data[ 2558] =  'sd74442;
    data[ 2559] =  'sd29571;
    data[ 2560] =  'sd43156;
    data[ 2561] = -'sd25590;
    data[ 2562] = -'sd15289;
    data[ 2563] =  'sd56818;
    data[ 2564] =  'sd70044;
    data[ 2565] = -'sd1215;
    data[ 2566] = -'sd8505;
    data[ 2567] = -'sd59535;
    data[ 2568] =  'sd74778;
    data[ 2569] =  'sd31923;
    data[ 2570] =  'sd59620;
    data[ 2571] = -'sd74183;
    data[ 2572] = -'sd27758;
    data[ 2573] = -'sd30465;
    data[ 2574] = -'sd49414;
    data[ 2575] = -'sd18216;
    data[ 2576] =  'sd36329;
    data[ 2577] = -'sd73379;
    data[ 2578] = -'sd22130;
    data[ 2579] =  'sd8931;
    data[ 2580] =  'sd62517;
    data[ 2581] = -'sd53904;
    data[ 2582] = -'sd49646;
    data[ 2583] = -'sd19840;
    data[ 2584] =  'sd24961;
    data[ 2585] =  'sd10886;
    data[ 2586] =  'sd76202;
    data[ 2587] =  'sd41891;
    data[ 2588] = -'sd34445;
    data[ 2589] = -'sd77274;
    data[ 2590] = -'sd49395;
    data[ 2591] = -'sd18083;
    data[ 2592] =  'sd37260;
    data[ 2593] = -'sd66862;
    data[ 2594] =  'sd23489;
    data[ 2595] =  'sd582;
    data[ 2596] =  'sd4074;
    data[ 2597] =  'sd28518;
    data[ 2598] =  'sd35785;
    data[ 2599] = -'sd77187;
    data[ 2600] = -'sd48786;
    data[ 2601] = -'sd13820;
    data[ 2602] =  'sd67101;
    data[ 2603] = -'sd21816;
    data[ 2604] =  'sd11129;
    data[ 2605] =  'sd77903;
    data[ 2606] =  'sd53798;
    data[ 2607] =  'sd48904;
    data[ 2608] =  'sd14646;
    data[ 2609] = -'sd61319;
    data[ 2610] =  'sd62290;
    data[ 2611] = -'sd55493;
    data[ 2612] = -'sd60769;
    data[ 2613] =  'sd66140;
    data[ 2614] = -'sd28543;
    data[ 2615] = -'sd35960;
    data[ 2616] =  'sd75962;
    data[ 2617] =  'sd40211;
    data[ 2618] = -'sd46205;
    data[ 2619] =  'sd4247;
    data[ 2620] =  'sd29729;
    data[ 2621] =  'sd44262;
    data[ 2622] = -'sd17848;
    data[ 2623] =  'sd38905;
    data[ 2624] = -'sd55347;
    data[ 2625] = -'sd59747;
    data[ 2626] =  'sd73294;
    data[ 2627] =  'sd21535;
    data[ 2628] = -'sd13096;
    data[ 2629] =  'sd72169;
    data[ 2630] =  'sd13660;
    data[ 2631] = -'sd68221;
    data[ 2632] =  'sd13976;
    data[ 2633] = -'sd66009;
    data[ 2634] =  'sd29460;
    data[ 2635] =  'sd42379;
    data[ 2636] = -'sd31029;
    data[ 2637] = -'sd53362;
    data[ 2638] = -'sd45852;
    data[ 2639] =  'sd6718;
    data[ 2640] =  'sd47026;
    data[ 2641] =  'sd1500;
    data[ 2642] =  'sd10500;
    data[ 2643] =  'sd73500;
    data[ 2644] =  'sd22977;
    data[ 2645] = -'sd3002;
    data[ 2646] = -'sd21014;
    data[ 2647] =  'sd16743;
    data[ 2648] = -'sd46640;
    data[ 2649] =  'sd1202;
    data[ 2650] =  'sd8414;
    data[ 2651] =  'sd58898;
    data[ 2652] = -'sd79237;
    data[ 2653] = -'sd63136;
    data[ 2654] =  'sd49571;
    data[ 2655] =  'sd19315;
    data[ 2656] = -'sd28636;
    data[ 2657] = -'sd36611;
    data[ 2658] =  'sd71405;
    data[ 2659] =  'sd8312;
    data[ 2660] =  'sd58184;
    data[ 2661] =  'sd79606;
    data[ 2662] =  'sd65719;
    data[ 2663] = -'sd31490;
    data[ 2664] = -'sd56589;
    data[ 2665] = -'sd68441;
    data[ 2666] =  'sd12436;
    data[ 2667] = -'sd76789;
    data[ 2668] = -'sd46000;
    data[ 2669] =  'sd5682;
    data[ 2670] =  'sd39774;
    data[ 2671] = -'sd49264;
    data[ 2672] = -'sd17166;
    data[ 2673] =  'sd43679;
    data[ 2674] = -'sd21929;
    data[ 2675] =  'sd10338;
    data[ 2676] =  'sd72366;
    data[ 2677] =  'sd15039;
    data[ 2678] = -'sd58568;
    data[ 2679] =  'sd81547;
    data[ 2680] =  'sd79306;
    data[ 2681] =  'sd63619;
    data[ 2682] = -'sd46190;
    data[ 2683] =  'sd4352;
    data[ 2684] =  'sd30464;
    data[ 2685] =  'sd49407;
    data[ 2686] =  'sd18167;
    data[ 2687] = -'sd36672;
    data[ 2688] =  'sd70978;
    data[ 2689] =  'sd5323;
    data[ 2690] =  'sd37261;
    data[ 2691] = -'sd66855;
    data[ 2692] =  'sd23538;
    data[ 2693] =  'sd925;
    data[ 2694] =  'sd6475;
    data[ 2695] =  'sd45325;
    data[ 2696] = -'sd10407;
    data[ 2697] = -'sd72849;
    data[ 2698] = -'sd18420;
    data[ 2699] =  'sd34901;
    data[ 2700] =  'sd80466;
    data[ 2701] =  'sd71739;
    data[ 2702] =  'sd10650;
    data[ 2703] =  'sd74550;
    data[ 2704] =  'sd30327;
    data[ 2705] =  'sd48448;
    data[ 2706] =  'sd11454;
    data[ 2707] =  'sd80178;
    data[ 2708] =  'sd69723;
    data[ 2709] = -'sd3462;
    data[ 2710] = -'sd24234;
    data[ 2711] = -'sd5797;
    data[ 2712] = -'sd40579;
    data[ 2713] =  'sd43629;
    data[ 2714] = -'sd22279;
    data[ 2715] =  'sd7888;
    data[ 2716] =  'sd55216;
    data[ 2717] =  'sd58830;
    data[ 2718] = -'sd79713;
    data[ 2719] = -'sd66468;
    data[ 2720] =  'sd26247;
    data[ 2721] =  'sd19888;
    data[ 2722] = -'sd24625;
    data[ 2723] = -'sd8534;
    data[ 2724] = -'sd59738;
    data[ 2725] =  'sd73357;
    data[ 2726] =  'sd21976;
    data[ 2727] = -'sd10009;
    data[ 2728] = -'sd70063;
    data[ 2729] =  'sd1082;
    data[ 2730] =  'sd7574;
    data[ 2731] =  'sd53018;
    data[ 2732] =  'sd43444;
    data[ 2733] = -'sd23574;
    data[ 2734] = -'sd1177;
    data[ 2735] = -'sd8239;
    data[ 2736] = -'sd57673;
    data[ 2737] = -'sd76029;
    data[ 2738] = -'sd40680;
    data[ 2739] =  'sd42922;
    data[ 2740] = -'sd27228;
    data[ 2741] = -'sd26755;
    data[ 2742] = -'sd23444;
    data[ 2743] = -'sd267;
    data[ 2744] = -'sd1869;
    data[ 2745] = -'sd13083;
    data[ 2746] =  'sd72260;
    data[ 2747] =  'sd14297;
    data[ 2748] = -'sd63762;
    data[ 2749] =  'sd45189;
    data[ 2750] = -'sd11359;
    data[ 2751] = -'sd79513;
    data[ 2752] = -'sd65068;
    data[ 2753] =  'sd36047;
    data[ 2754] = -'sd75353;
    data[ 2755] = -'sd35948;
    data[ 2756] =  'sd76046;
    data[ 2757] =  'sd40799;
    data[ 2758] = -'sd42089;
    data[ 2759] =  'sd33059;
    data[ 2760] =  'sd67572;
    data[ 2761] = -'sd18519;
    data[ 2762] =  'sd34208;
    data[ 2763] =  'sd75615;
    data[ 2764] =  'sd37782;
    data[ 2765] = -'sd63208;
    data[ 2766] =  'sd49067;
    data[ 2767] =  'sd15787;
    data[ 2768] = -'sd53332;
    data[ 2769] = -'sd45642;
    data[ 2770] =  'sd8188;
    data[ 2771] =  'sd57316;
    data[ 2772] =  'sd73530;
    data[ 2773] =  'sd23187;
    data[ 2774] = -'sd1532;
    data[ 2775] = -'sd10724;
    data[ 2776] = -'sd75068;
    data[ 2777] = -'sd33953;
    data[ 2778] = -'sd73830;
    data[ 2779] = -'sd25287;
    data[ 2780] = -'sd13168;
    data[ 2781] =  'sd71665;
    data[ 2782] =  'sd10132;
    data[ 2783] =  'sd70924;
    data[ 2784] =  'sd4945;
    data[ 2785] =  'sd34615;
    data[ 2786] =  'sd78464;
    data[ 2787] =  'sd57725;
    data[ 2788] =  'sd76393;
    data[ 2789] =  'sd43228;
    data[ 2790] = -'sd25086;
    data[ 2791] = -'sd11761;
    data[ 2792] =  'sd81514;
    data[ 2793] =  'sd79075;
    data[ 2794] =  'sd62002;
    data[ 2795] = -'sd57509;
    data[ 2796] = -'sd74881;
    data[ 2797] = -'sd32644;
    data[ 2798] = -'sd64667;
    data[ 2799] =  'sd38854;
    data[ 2800] = -'sd55704;
    data[ 2801] = -'sd62246;
    data[ 2802] =  'sd55801;
    data[ 2803] =  'sd62925;
    data[ 2804] = -'sd51048;
    data[ 2805] = -'sd29654;
    data[ 2806] = -'sd43737;
    data[ 2807] =  'sd21523;
    data[ 2808] = -'sd13180;
    data[ 2809] =  'sd71581;
    data[ 2810] =  'sd9544;
    data[ 2811] =  'sd66808;
    data[ 2812] = -'sd23867;
    data[ 2813] = -'sd3228;
    data[ 2814] = -'sd22596;
    data[ 2815] =  'sd5669;
    data[ 2816] =  'sd39683;
    data[ 2817] = -'sd49901;
    data[ 2818] = -'sd21625;
    data[ 2819] =  'sd12466;
    data[ 2820] = -'sd76579;
    data[ 2821] = -'sd44530;
    data[ 2822] =  'sd15972;
    data[ 2823] = -'sd52037;
    data[ 2824] = -'sd36577;
    data[ 2825] =  'sd71643;
    data[ 2826] =  'sd9978;
    data[ 2827] =  'sd69846;
    data[ 2828] = -'sd2601;
    data[ 2829] = -'sd18207;
    data[ 2830] =  'sd36392;
    data[ 2831] = -'sd72938;
    data[ 2832] = -'sd19043;
    data[ 2833] =  'sd30540;
    data[ 2834] =  'sd49939;
    data[ 2835] =  'sd21891;
    data[ 2836] = -'sd10604;
    data[ 2837] = -'sd74228;
    data[ 2838] = -'sd28073;
    data[ 2839] = -'sd32670;
    data[ 2840] = -'sd64849;
    data[ 2841] =  'sd37580;
    data[ 2842] = -'sd64622;
    data[ 2843] =  'sd39169;
    data[ 2844] = -'sd53499;
    data[ 2845] = -'sd46811;
    data[ 2846] =  'sd5;
    data[ 2847] =  'sd35;
    data[ 2848] =  'sd245;
    data[ 2849] =  'sd1715;
    data[ 2850] =  'sd12005;
    data[ 2851] = -'sd79806;
    data[ 2852] = -'sd67119;
    data[ 2853] =  'sd21690;
    data[ 2854] = -'sd12011;
    data[ 2855] =  'sd79764;
    data[ 2856] =  'sd66825;
    data[ 2857] = -'sd23748;
    data[ 2858] = -'sd2395;
    data[ 2859] = -'sd16765;
    data[ 2860] =  'sd46486;
    data[ 2861] = -'sd2280;
    data[ 2862] = -'sd15960;
    data[ 2863] =  'sd52121;
    data[ 2864] =  'sd37165;
    data[ 2865] = -'sd67527;
    data[ 2866] =  'sd18834;
    data[ 2867] = -'sd32003;
    data[ 2868] = -'sd60180;
    data[ 2869] =  'sd70263;
    data[ 2870] =  'sd318;
    data[ 2871] =  'sd2226;
    data[ 2872] =  'sd15582;
    data[ 2873] = -'sd54767;
    data[ 2874] = -'sd55687;
    data[ 2875] = -'sd62127;
    data[ 2876] =  'sd56634;
    data[ 2877] =  'sd68756;
    data[ 2878] = -'sd10231;
    data[ 2879] = -'sd71617;
    data[ 2880] = -'sd9796;
    data[ 2881] = -'sd68572;
    data[ 2882] =  'sd11519;
    data[ 2883] =  'sd80633;
    data[ 2884] =  'sd72908;
    data[ 2885] =  'sd18833;
    data[ 2886] = -'sd32010;
    data[ 2887] = -'sd60229;
    data[ 2888] =  'sd69920;
    data[ 2889] = -'sd2083;
    data[ 2890] = -'sd14581;
    data[ 2891] =  'sd61774;
    data[ 2892] = -'sd59105;
    data[ 2893] =  'sd77788;
    data[ 2894] =  'sd52993;
    data[ 2895] =  'sd43269;
    data[ 2896] = -'sd24799;
    data[ 2897] = -'sd9752;
    data[ 2898] = -'sd68264;
    data[ 2899] =  'sd13675;
    data[ 2900] = -'sd68116;
    data[ 2901] =  'sd14711;
    data[ 2902] = -'sd60864;
    data[ 2903] =  'sd65475;
    data[ 2904] = -'sd33198;
    data[ 2905] = -'sd68545;
    data[ 2906] =  'sd11708;
    data[ 2907] = -'sd81885;
    data[ 2908] = -'sd81672;
    data[ 2909] = -'sd80181;
    data[ 2910] = -'sd69744;
    data[ 2911] =  'sd3315;
    data[ 2912] =  'sd23205;
    data[ 2913] = -'sd1406;
    data[ 2914] = -'sd9842;
    data[ 2915] = -'sd68894;
    data[ 2916] =  'sd9265;
    data[ 2917] =  'sd64855;
    data[ 2918] = -'sd37538;
    data[ 2919] =  'sd64916;
    data[ 2920] = -'sd37111;
    data[ 2921] =  'sd67905;
    data[ 2922] = -'sd16188;
    data[ 2923] =  'sd50525;
    data[ 2924] =  'sd25993;
    data[ 2925] =  'sd18110;
    data[ 2926] = -'sd37071;
    data[ 2927] =  'sd68185;
    data[ 2928] = -'sd14228;
    data[ 2929] =  'sd64245;
    data[ 2930] = -'sd41808;
    data[ 2931] =  'sd35026;
    data[ 2932] =  'sd81341;
    data[ 2933] =  'sd77864;
    data[ 2934] =  'sd53525;
    data[ 2935] =  'sd46993;
    data[ 2936] =  'sd1269;
    data[ 2937] =  'sd8883;
    data[ 2938] =  'sd62181;
    data[ 2939] = -'sd56256;
    data[ 2940] = -'sd66110;
    data[ 2941] =  'sd28753;
    data[ 2942] =  'sd37430;
    data[ 2943] = -'sd65672;
    data[ 2944] =  'sd31819;
    data[ 2945] =  'sd58892;
    data[ 2946] = -'sd79279;
    data[ 2947] = -'sd63430;
    data[ 2948] =  'sd47513;
    data[ 2949] =  'sd4909;
    data[ 2950] =  'sd34363;
    data[ 2951] =  'sd76700;
    data[ 2952] =  'sd45377;
    data[ 2953] = -'sd10043;
    data[ 2954] = -'sd70301;
    data[ 2955] = -'sd584;
    data[ 2956] = -'sd4088;
    data[ 2957] = -'sd28616;
    data[ 2958] = -'sd36471;
    data[ 2959] =  'sd72385;
    data[ 2960] =  'sd15172;
    data[ 2961] = -'sd57637;
    data[ 2962] = -'sd75777;
    data[ 2963] = -'sd38916;
    data[ 2964] =  'sd55270;
    data[ 2965] =  'sd59208;
    data[ 2966] = -'sd77067;
    data[ 2967] = -'sd47946;
    data[ 2968] = -'sd7940;
    data[ 2969] = -'sd55580;
    data[ 2970] = -'sd61378;
    data[ 2971] =  'sd61877;
    data[ 2972] = -'sd58384;
    data[ 2973] = -'sd81006;
    data[ 2974] = -'sd75519;
    data[ 2975] = -'sd37110;
    data[ 2976] =  'sd67912;
    data[ 2977] = -'sd16139;
    data[ 2978] =  'sd50868;
    data[ 2979] =  'sd28394;
    data[ 2980] =  'sd34917;
    data[ 2981] =  'sd80578;
    data[ 2982] =  'sd72523;
    data[ 2983] =  'sd16138;
    data[ 2984] = -'sd50875;
    data[ 2985] = -'sd28443;
    data[ 2986] = -'sd35260;
    data[ 2987] =  'sd80862;
    data[ 2988] =  'sd74511;
    data[ 2989] =  'sd30054;
    data[ 2990] =  'sd46537;
    data[ 2991] = -'sd1923;
    data[ 2992] = -'sd13461;
    data[ 2993] =  'sd69614;
    data[ 2994] = -'sd4225;
    data[ 2995] = -'sd29575;
    data[ 2996] = -'sd43184;
    data[ 2997] =  'sd25394;
    data[ 2998] =  'sd13917;
    data[ 2999] = -'sd66422;
    data[ 3000] =  'sd26569;
    data[ 3001] =  'sd22142;
    data[ 3002] = -'sd8847;
    data[ 3003] = -'sd61929;
    data[ 3004] =  'sd58020;
    data[ 3005] =  'sd78458;
    data[ 3006] =  'sd57683;
    data[ 3007] =  'sd76099;
    data[ 3008] =  'sd41170;
    data[ 3009] = -'sd39492;
    data[ 3010] =  'sd51238;
    data[ 3011] =  'sd30984;
    data[ 3012] =  'sd53047;
    data[ 3013] =  'sd43647;
    data[ 3014] = -'sd22153;
    data[ 3015] =  'sd8770;
    data[ 3016] =  'sd61390;
    data[ 3017] = -'sd61793;
    data[ 3018] =  'sd58972;
    data[ 3019] = -'sd78719;
    data[ 3020] = -'sd59510;
    data[ 3021] =  'sd74953;
    data[ 3022] =  'sd33148;
    data[ 3023] =  'sd68195;
    data[ 3024] = -'sd14158;
    data[ 3025] =  'sd64735;
    data[ 3026] = -'sd38378;
    data[ 3027] =  'sd59036;
    data[ 3028] = -'sd78271;
    data[ 3029] = -'sd56374;
    data[ 3030] = -'sd66936;
    data[ 3031] =  'sd22971;
    data[ 3032] = -'sd3044;
    data[ 3033] = -'sd21308;
    data[ 3034] =  'sd14685;
    data[ 3035] = -'sd61046;
    data[ 3036] =  'sd64201;
    data[ 3037] = -'sd42116;
    data[ 3038] =  'sd32870;
    data[ 3039] =  'sd66249;
    data[ 3040] = -'sd27780;
    data[ 3041] = -'sd30619;
    data[ 3042] = -'sd50492;
    data[ 3043] = -'sd25762;
    data[ 3044] = -'sd16493;
    data[ 3045] =  'sd48390;
    data[ 3046] =  'sd11048;
    data[ 3047] =  'sd77336;
    data[ 3048] =  'sd49829;
    data[ 3049] =  'sd21121;
    data[ 3050] = -'sd15994;
    data[ 3051] =  'sd51883;
    data[ 3052] =  'sd35499;
    data[ 3053] = -'sd79189;
    data[ 3054] = -'sd62800;
    data[ 3055] =  'sd51923;
    data[ 3056] =  'sd35779;
    data[ 3057] = -'sd77229;
    data[ 3058] = -'sd49080;
    data[ 3059] = -'sd15878;
    data[ 3060] =  'sd52695;
    data[ 3061] =  'sd41183;
    data[ 3062] = -'sd39401;
    data[ 3063] =  'sd51875;
    data[ 3064] =  'sd35443;
    data[ 3065] = -'sd79581;
    data[ 3066] = -'sd65544;
    data[ 3067] =  'sd32715;
    data[ 3068] =  'sd65164;
    data[ 3069] = -'sd35375;
    data[ 3070] =  'sd80057;
    data[ 3071] =  'sd68876;
    data[ 3072] = -'sd9391;
    data[ 3073] = -'sd65737;
    data[ 3074] =  'sd31364;
    data[ 3075] =  'sd55707;
    data[ 3076] =  'sd62267;
    data[ 3077] = -'sd55654;
    data[ 3078] = -'sd61896;
    data[ 3079] =  'sd58251;
    data[ 3080] =  'sd80075;
    data[ 3081] =  'sd69002;
    data[ 3082] = -'sd8509;
    data[ 3083] = -'sd59563;
    data[ 3084] =  'sd74582;
    data[ 3085] =  'sd30551;
    data[ 3086] =  'sd50016;
    data[ 3087] =  'sd22430;
    data[ 3088] = -'sd6831;
    data[ 3089] = -'sd47817;
    data[ 3090] = -'sd7037;
    data[ 3091] = -'sd49259;
    data[ 3092] = -'sd17131;
    data[ 3093] =  'sd43924;
    data[ 3094] = -'sd20214;
    data[ 3095] =  'sd22343;
    data[ 3096] = -'sd7440;
    data[ 3097] = -'sd52080;
    data[ 3098] = -'sd36878;
    data[ 3099] =  'sd69536;
    data[ 3100] = -'sd4771;
    data[ 3101] = -'sd33397;
    data[ 3102] = -'sd69938;
    data[ 3103] =  'sd1957;
    data[ 3104] =  'sd13699;
    data[ 3105] = -'sd67948;
    data[ 3106] =  'sd15887;
    data[ 3107] = -'sd52632;
    data[ 3108] = -'sd40742;
    data[ 3109] =  'sd42488;
    data[ 3110] = -'sd30266;
    data[ 3111] = -'sd48021;
    data[ 3112] = -'sd8465;
    data[ 3113] = -'sd59255;
    data[ 3114] =  'sd76738;
    data[ 3115] =  'sd45643;
    data[ 3116] = -'sd8181;
    data[ 3117] = -'sd57267;
    data[ 3118] = -'sd73187;
    data[ 3119] = -'sd20786;
    data[ 3120] =  'sd18339;
    data[ 3121] = -'sd35468;
    data[ 3122] =  'sd79406;
    data[ 3123] =  'sd64319;
    data[ 3124] = -'sd41290;
    data[ 3125] =  'sd38652;
    data[ 3126] = -'sd57118;
    data[ 3127] = -'sd72144;
    data[ 3128] = -'sd13485;
    data[ 3129] =  'sd69446;
    data[ 3130] = -'sd5401;
    data[ 3131] = -'sd37807;
    data[ 3132] =  'sd63033;
    data[ 3133] = -'sd50292;
    data[ 3134] = -'sd24362;
    data[ 3135] = -'sd6693;
    data[ 3136] = -'sd46851;
    data[ 3137] = -'sd275;
    data[ 3138] = -'sd1925;
    data[ 3139] = -'sd13475;
    data[ 3140] =  'sd69516;
    data[ 3141] = -'sd4911;
    data[ 3142] = -'sd34377;
    data[ 3143] = -'sd76798;
    data[ 3144] = -'sd46063;
    data[ 3145] =  'sd5241;
    data[ 3146] =  'sd36687;
    data[ 3147] = -'sd70873;
    data[ 3148] = -'sd4588;
    data[ 3149] = -'sd32116;
    data[ 3150] = -'sd60971;
    data[ 3151] =  'sd64726;
    data[ 3152] = -'sd38441;
    data[ 3153] =  'sd58595;
    data[ 3154] = -'sd81358;
    data[ 3155] = -'sd77983;
    data[ 3156] = -'sd54358;
    data[ 3157] = -'sd52824;
    data[ 3158] = -'sd42086;
    data[ 3159] =  'sd33080;
    data[ 3160] =  'sd67719;
    data[ 3161] = -'sd17490;
    data[ 3162] =  'sd41411;
    data[ 3163] = -'sd37805;
    data[ 3164] =  'sd63047;
    data[ 3165] = -'sd50194;
    data[ 3166] = -'sd23676;
    data[ 3167] = -'sd1891;
    data[ 3168] = -'sd13237;
    data[ 3169] =  'sd71182;
    data[ 3170] =  'sd6751;
    data[ 3171] =  'sd47257;
    data[ 3172] =  'sd3117;
    data[ 3173] =  'sd21819;
    data[ 3174] = -'sd11108;
    data[ 3175] = -'sd77756;
    data[ 3176] = -'sd52769;
    data[ 3177] = -'sd41701;
    data[ 3178] =  'sd35775;
    data[ 3179] = -'sd77257;
    data[ 3180] = -'sd49276;
    data[ 3181] = -'sd17250;
    data[ 3182] =  'sd43091;
    data[ 3183] = -'sd26045;
    data[ 3184] = -'sd18474;
    data[ 3185] =  'sd34523;
    data[ 3186] =  'sd77820;
    data[ 3187] =  'sd53217;
    data[ 3188] =  'sd44837;
    data[ 3189] = -'sd13823;
    data[ 3190] =  'sd67080;
    data[ 3191] = -'sd21963;
    data[ 3192] =  'sd10100;
    data[ 3193] =  'sd70700;
    data[ 3194] =  'sd3377;
    data[ 3195] =  'sd23639;
    data[ 3196] =  'sd1632;
    data[ 3197] =  'sd11424;
    data[ 3198] =  'sd79968;
    data[ 3199] =  'sd68253;
    data[ 3200] = -'sd13752;
    data[ 3201] =  'sd67577;
    data[ 3202] = -'sd18484;
    data[ 3203] =  'sd34453;
    data[ 3204] =  'sd77330;
    data[ 3205] =  'sd49787;
    data[ 3206] =  'sd20827;
    data[ 3207] = -'sd18052;
    data[ 3208] =  'sd37477;
    data[ 3209] = -'sd65343;
    data[ 3210] =  'sd34122;
    data[ 3211] =  'sd75013;
    data[ 3212] =  'sd33568;
    data[ 3213] =  'sd71135;
    data[ 3214] =  'sd6422;
    data[ 3215] =  'sd44954;
    data[ 3216] = -'sd13004;
    data[ 3217] =  'sd72813;
    data[ 3218] =  'sd18168;
    data[ 3219] = -'sd36665;
    data[ 3220] =  'sd71027;
    data[ 3221] =  'sd5666;
    data[ 3222] =  'sd39662;
    data[ 3223] = -'sd50048;
    data[ 3224] = -'sd22654;
    data[ 3225] =  'sd5263;
    data[ 3226] =  'sd36841;
    data[ 3227] = -'sd69795;
    data[ 3228] =  'sd2958;
    data[ 3229] =  'sd20706;
    data[ 3230] = -'sd18899;
    data[ 3231] =  'sd31548;
    data[ 3232] =  'sd56995;
    data[ 3233] =  'sd71283;
    data[ 3234] =  'sd7458;
    data[ 3235] =  'sd52206;
    data[ 3236] =  'sd37760;
    data[ 3237] = -'sd63362;
    data[ 3238] =  'sd47989;
    data[ 3239] =  'sd8241;
    data[ 3240] =  'sd57687;
    data[ 3241] =  'sd76127;
    data[ 3242] =  'sd41366;
    data[ 3243] = -'sd38120;
    data[ 3244] =  'sd60842;
    data[ 3245] = -'sd65629;
    data[ 3246] =  'sd32120;
    data[ 3247] =  'sd60999;
    data[ 3248] = -'sd64530;
    data[ 3249] =  'sd39813;
    data[ 3250] = -'sd48991;
    data[ 3251] = -'sd15255;
    data[ 3252] =  'sd57056;
    data[ 3253] =  'sd71710;
    data[ 3254] =  'sd10447;
    data[ 3255] =  'sd73129;
    data[ 3256] =  'sd20380;
    data[ 3257] = -'sd21181;
    data[ 3258] =  'sd15574;
    data[ 3259] = -'sd54823;
    data[ 3260] = -'sd56079;
    data[ 3261] = -'sd64871;
    data[ 3262] =  'sd37426;
    data[ 3263] = -'sd65700;
    data[ 3264] =  'sd31623;
    data[ 3265] =  'sd57520;
    data[ 3266] =  'sd74958;
    data[ 3267] =  'sd33183;
    data[ 3268] =  'sd68440;
    data[ 3269] = -'sd12443;
    data[ 3270] =  'sd76740;
    data[ 3271] =  'sd45657;
    data[ 3272] = -'sd8083;
    data[ 3273] = -'sd56581;
    data[ 3274] = -'sd68385;
    data[ 3275] =  'sd12828;
    data[ 3276] = -'sd74045;
    data[ 3277] = -'sd26792;
    data[ 3278] = -'sd23703;
    data[ 3279] = -'sd2080;
    data[ 3280] = -'sd14560;
    data[ 3281] =  'sd61921;
    data[ 3282] = -'sd58076;
    data[ 3283] = -'sd78850;
    data[ 3284] = -'sd60427;
    data[ 3285] =  'sd68534;
    data[ 3286] = -'sd11785;
    data[ 3287] =  'sd81346;
    data[ 3288] =  'sd77899;
    data[ 3289] =  'sd53770;
    data[ 3290] =  'sd48708;
    data[ 3291] =  'sd13274;
    data[ 3292] = -'sd70923;
    data[ 3293] = -'sd4938;
    data[ 3294] = -'sd34566;
    data[ 3295] = -'sd78121;
    data[ 3296] = -'sd55324;
    data[ 3297] = -'sd59586;
    data[ 3298] =  'sd74421;
    data[ 3299] =  'sd29424;
    data[ 3300] =  'sd42127;
    data[ 3301] = -'sd32793;
    data[ 3302] = -'sd65710;
    data[ 3303] =  'sd31553;
    data[ 3304] =  'sd57030;
    data[ 3305] =  'sd71528;
    data[ 3306] =  'sd9173;
    data[ 3307] =  'sd64211;
    data[ 3308] = -'sd42046;
    data[ 3309] =  'sd33360;
    data[ 3310] =  'sd69679;
    data[ 3311] = -'sd3770;
    data[ 3312] = -'sd26390;
    data[ 3313] = -'sd20889;
    data[ 3314] =  'sd17618;
    data[ 3315] = -'sd40515;
    data[ 3316] =  'sd44077;
    data[ 3317] = -'sd19143;
    data[ 3318] =  'sd29840;
    data[ 3319] =  'sd45039;
    data[ 3320] = -'sd12409;
    data[ 3321] =  'sd76978;
    data[ 3322] =  'sd47323;
    data[ 3323] =  'sd3579;
    data[ 3324] =  'sd25053;
    data[ 3325] =  'sd11530;
    data[ 3326] =  'sd80710;
    data[ 3327] =  'sd73447;
    data[ 3328] =  'sd22606;
    data[ 3329] = -'sd5599;
    data[ 3330] = -'sd39193;
    data[ 3331] =  'sd53331;
    data[ 3332] =  'sd45635;
    data[ 3333] = -'sd8237;
    data[ 3334] = -'sd57659;
    data[ 3335] = -'sd75931;
    data[ 3336] = -'sd39994;
    data[ 3337] =  'sd47724;
    data[ 3338] =  'sd6386;
    data[ 3339] =  'sd44702;
    data[ 3340] = -'sd14768;
    data[ 3341] =  'sd60465;
    data[ 3342] = -'sd68268;
    data[ 3343] =  'sd13647;
    data[ 3344] = -'sd68312;
    data[ 3345] =  'sd13339;
    data[ 3346] = -'sd70468;
    data[ 3347] = -'sd1753;
    data[ 3348] = -'sd12271;
    data[ 3349] =  'sd77944;
    data[ 3350] =  'sd54085;
    data[ 3351] =  'sd50913;
    data[ 3352] =  'sd28709;
    data[ 3353] =  'sd37122;
    data[ 3354] = -'sd67828;
    data[ 3355] =  'sd16727;
    data[ 3356] = -'sd46752;
    data[ 3357] =  'sd418;
    data[ 3358] =  'sd2926;
    data[ 3359] =  'sd20482;
    data[ 3360] = -'sd20467;
    data[ 3361] =  'sd20572;
    data[ 3362] = -'sd19837;
    data[ 3363] =  'sd24982;
    data[ 3364] =  'sd11033;
    data[ 3365] =  'sd77231;
    data[ 3366] =  'sd49094;
    data[ 3367] =  'sd15976;
    data[ 3368] = -'sd52009;
    data[ 3369] = -'sd36381;
    data[ 3370] =  'sd73015;
    data[ 3371] =  'sd19582;
    data[ 3372] = -'sd26767;
    data[ 3373] = -'sd23528;
    data[ 3374] = -'sd855;
    data[ 3375] = -'sd5985;
    data[ 3376] = -'sd41895;
    data[ 3377] =  'sd34417;
    data[ 3378] =  'sd77078;
    data[ 3379] =  'sd48023;
    data[ 3380] =  'sd8479;
    data[ 3381] =  'sd59353;
    data[ 3382] = -'sd76052;
    data[ 3383] = -'sd40841;
    data[ 3384] =  'sd41795;
    data[ 3385] = -'sd35117;
    data[ 3386] =  'sd81863;
    data[ 3387] =  'sd81518;
    data[ 3388] =  'sd79103;
    data[ 3389] =  'sd62198;
    data[ 3390] = -'sd56137;
    data[ 3391] = -'sd65277;
    data[ 3392] =  'sd34584;
    data[ 3393] =  'sd78247;
    data[ 3394] =  'sd56206;
    data[ 3395] =  'sd65760;
    data[ 3396] = -'sd31203;
    data[ 3397] = -'sd54580;
    data[ 3398] = -'sd54378;
    data[ 3399] = -'sd52964;
    data[ 3400] = -'sd43066;
    data[ 3401] =  'sd26220;
    data[ 3402] =  'sd19699;
    data[ 3403] = -'sd25948;
    data[ 3404] = -'sd17795;
    data[ 3405] =  'sd39276;
    data[ 3406] = -'sd52750;
    data[ 3407] = -'sd41568;
    data[ 3408] =  'sd36706;
    data[ 3409] = -'sd70740;
    data[ 3410] = -'sd3657;
    data[ 3411] = -'sd25599;
    data[ 3412] = -'sd15352;
    data[ 3413] =  'sd56377;
    data[ 3414] =  'sd66957;
    data[ 3415] = -'sd22824;
    data[ 3416] =  'sd4073;
    data[ 3417] =  'sd28511;
    data[ 3418] =  'sd35736;
    data[ 3419] = -'sd77530;
    data[ 3420] = -'sd51187;
    data[ 3421] = -'sd30627;
    data[ 3422] = -'sd50548;
    data[ 3423] = -'sd26154;
    data[ 3424] = -'sd19237;
    data[ 3425] =  'sd29182;
    data[ 3426] =  'sd40433;
    data[ 3427] = -'sd44651;
    data[ 3428] =  'sd15125;
    data[ 3429] = -'sd57966;
    data[ 3430] = -'sd78080;
    data[ 3431] = -'sd55037;
    data[ 3432] = -'sd57577;
    data[ 3433] = -'sd75357;
    data[ 3434] = -'sd35976;
    data[ 3435] =  'sd75850;
    data[ 3436] =  'sd39427;
    data[ 3437] = -'sd51693;
    data[ 3438] = -'sd34169;
    data[ 3439] = -'sd75342;
    data[ 3440] = -'sd35871;
    data[ 3441] =  'sd76585;
    data[ 3442] =  'sd44572;
    data[ 3443] = -'sd15678;
    data[ 3444] =  'sd54095;
    data[ 3445] =  'sd50983;
    data[ 3446] =  'sd29199;
    data[ 3447] =  'sd40552;
    data[ 3448] = -'sd43818;
    data[ 3449] =  'sd20956;
    data[ 3450] = -'sd17149;
    data[ 3451] =  'sd43798;
    data[ 3452] = -'sd21096;
    data[ 3453] =  'sd16169;
    data[ 3454] = -'sd50658;
    data[ 3455] = -'sd26924;
    data[ 3456] = -'sd24627;
    data[ 3457] = -'sd8548;
    data[ 3458] = -'sd59836;
    data[ 3459] =  'sd72671;
    data[ 3460] =  'sd17174;
    data[ 3461] = -'sd43623;
    data[ 3462] =  'sd22321;
    data[ 3463] = -'sd7594;
    data[ 3464] = -'sd53158;
    data[ 3465] = -'sd44424;
    data[ 3466] =  'sd16714;
    data[ 3467] = -'sd46843;
    data[ 3468] = -'sd219;
    data[ 3469] = -'sd1533;
    data[ 3470] = -'sd10731;
    data[ 3471] = -'sd75117;
    data[ 3472] = -'sd34296;
    data[ 3473] = -'sd76231;
    data[ 3474] = -'sd42094;
    data[ 3475] =  'sd33024;
    data[ 3476] =  'sd67327;
    data[ 3477] = -'sd20234;
    data[ 3478] =  'sd22203;
    data[ 3479] = -'sd8420;
    data[ 3480] = -'sd58940;
    data[ 3481] =  'sd78943;
    data[ 3482] =  'sd61078;
    data[ 3483] = -'sd63977;
    data[ 3484] =  'sd43684;
    data[ 3485] = -'sd21894;
    data[ 3486] =  'sd10583;
    data[ 3487] =  'sd74081;
    data[ 3488] =  'sd27044;
    data[ 3489] =  'sd25467;
    data[ 3490] =  'sd14428;
    data[ 3491] = -'sd62845;
    data[ 3492] =  'sd51608;
    data[ 3493] =  'sd33574;
    data[ 3494] =  'sd71177;
    data[ 3495] =  'sd6716;
    data[ 3496] =  'sd47012;
    data[ 3497] =  'sd1402;
    data[ 3498] =  'sd9814;
    data[ 3499] =  'sd68698;
    data[ 3500] = -'sd10637;
    data[ 3501] = -'sd74459;
    data[ 3502] = -'sd29690;
    data[ 3503] = -'sd43989;
    data[ 3504] =  'sd19759;
    data[ 3505] = -'sd25528;
    data[ 3506] = -'sd14855;
    data[ 3507] =  'sd59856;
    data[ 3508] = -'sd72531;
    data[ 3509] = -'sd16194;
    data[ 3510] =  'sd50483;
    data[ 3511] =  'sd25699;
    data[ 3512] =  'sd16052;
    data[ 3513] = -'sd51477;
    data[ 3514] = -'sd32657;
    data[ 3515] = -'sd64758;
    data[ 3516] =  'sd38217;
    data[ 3517] = -'sd60163;
    data[ 3518] =  'sd70382;
    data[ 3519] =  'sd1151;
    data[ 3520] =  'sd8057;
    data[ 3521] =  'sd56399;
    data[ 3522] =  'sd67111;
    data[ 3523] = -'sd21746;
    data[ 3524] =  'sd11619;
    data[ 3525] =  'sd81333;
    data[ 3526] =  'sd77808;
    data[ 3527] =  'sd53133;
    data[ 3528] =  'sd44249;
    data[ 3529] = -'sd17939;
    data[ 3530] =  'sd38268;
    data[ 3531] = -'sd59806;
    data[ 3532] =  'sd72881;
    data[ 3533] =  'sd18644;
    data[ 3534] = -'sd33333;
    data[ 3535] = -'sd69490;
    data[ 3536] =  'sd5093;
    data[ 3537] =  'sd35651;
    data[ 3538] = -'sd78125;
    data[ 3539] = -'sd55352;
    data[ 3540] = -'sd59782;
    data[ 3541] =  'sd73049;
    data[ 3542] =  'sd19820;
    data[ 3543] = -'sd25101;
    data[ 3544] = -'sd11866;
    data[ 3545] =  'sd80779;
    data[ 3546] =  'sd73930;
    data[ 3547] =  'sd25987;
    data[ 3548] =  'sd18068;
    data[ 3549] = -'sd37365;
    data[ 3550] =  'sd66127;
    data[ 3551] = -'sd28634;
    data[ 3552] = -'sd36597;
    data[ 3553] =  'sd71503;
    data[ 3554] =  'sd8998;
    data[ 3555] =  'sd62986;
    data[ 3556] = -'sd50621;
    data[ 3557] = -'sd26665;
    data[ 3558] = -'sd22814;
    data[ 3559] =  'sd4143;
    data[ 3560] =  'sd29001;
    data[ 3561] =  'sd39166;
    data[ 3562] = -'sd53520;
    data[ 3563] = -'sd46958;
    data[ 3564] = -'sd1024;
    data[ 3565] = -'sd7168;
    data[ 3566] = -'sd50176;
    data[ 3567] = -'sd23550;
    data[ 3568] = -'sd1009;
    data[ 3569] = -'sd7063;
    data[ 3570] = -'sd49441;
    data[ 3571] = -'sd18405;
    data[ 3572] =  'sd35006;
    data[ 3573] =  'sd81201;
    data[ 3574] =  'sd76884;
    data[ 3575] =  'sd46665;
    data[ 3576] = -'sd1027;
    data[ 3577] = -'sd7189;
    data[ 3578] = -'sd50323;
    data[ 3579] = -'sd24579;
    data[ 3580] = -'sd8212;
    data[ 3581] = -'sd57484;
    data[ 3582] = -'sd74706;
    data[ 3583] = -'sd31419;
    data[ 3584] = -'sd56092;
    data[ 3585] = -'sd64962;
    data[ 3586] =  'sd36789;
    data[ 3587] = -'sd70159;
    data[ 3588] =  'sd410;
    data[ 3589] =  'sd2870;
    data[ 3590] =  'sd20090;
    data[ 3591] = -'sd23211;
    data[ 3592] =  'sd1364;
    data[ 3593] =  'sd9548;
    data[ 3594] =  'sd66836;
    data[ 3595] = -'sd23671;
    data[ 3596] = -'sd1856;
    data[ 3597] = -'sd12992;
    data[ 3598] =  'sd72897;
    data[ 3599] =  'sd18756;
    data[ 3600] = -'sd32549;
    data[ 3601] = -'sd64002;
    data[ 3602] =  'sd43509;
    data[ 3603] = -'sd23119;
    data[ 3604] =  'sd2008;
    data[ 3605] =  'sd14056;
    data[ 3606] = -'sd65449;
    data[ 3607] =  'sd33380;
    data[ 3608] =  'sd69819;
    data[ 3609] = -'sd2790;
    data[ 3610] = -'sd19530;
    data[ 3611] =  'sd27131;
    data[ 3612] =  'sd26076;
    data[ 3613] =  'sd18691;
    data[ 3614] = -'sd33004;
    data[ 3615] = -'sd67187;
    data[ 3616] =  'sd21214;
    data[ 3617] = -'sd15343;
    data[ 3618] =  'sd56440;
    data[ 3619] =  'sd67398;
    data[ 3620] = -'sd19737;
    data[ 3621] =  'sd25682;
    data[ 3622] =  'sd15933;
    data[ 3623] = -'sd52310;
    data[ 3624] = -'sd38488;
    data[ 3625] =  'sd58266;
    data[ 3626] =  'sd80180;
    data[ 3627] =  'sd69737;
    data[ 3628] = -'sd3364;
    data[ 3629] = -'sd23548;
    data[ 3630] = -'sd995;
    data[ 3631] = -'sd6965;
    data[ 3632] = -'sd48755;
    data[ 3633] = -'sd13603;
    data[ 3634] =  'sd68620;
    data[ 3635] = -'sd11183;
    data[ 3636] = -'sd78281;
    data[ 3637] = -'sd56444;
    data[ 3638] = -'sd67426;
    data[ 3639] =  'sd19541;
    data[ 3640] = -'sd27054;
    data[ 3641] = -'sd25537;
    data[ 3642] = -'sd14918;
    data[ 3643] =  'sd59415;
    data[ 3644] = -'sd75618;
    data[ 3645] = -'sd37803;
    data[ 3646] =  'sd63061;
    data[ 3647] = -'sd50096;
    data[ 3648] = -'sd22990;
    data[ 3649] =  'sd2911;
    data[ 3650] =  'sd20377;
    data[ 3651] = -'sd21202;
    data[ 3652] =  'sd15427;
    data[ 3653] = -'sd55852;
    data[ 3654] = -'sd63282;
    data[ 3655] =  'sd48549;
    data[ 3656] =  'sd12161;
    data[ 3657] = -'sd78714;
    data[ 3658] = -'sd59475;
    data[ 3659] =  'sd75198;
    data[ 3660] =  'sd34863;
    data[ 3661] =  'sd80200;
    data[ 3662] =  'sd69877;
    data[ 3663] = -'sd2384;
    data[ 3664] = -'sd16688;
    data[ 3665] =  'sd47025;
    data[ 3666] =  'sd1493;
    data[ 3667] =  'sd10451;
    data[ 3668] =  'sd73157;
    data[ 3669] =  'sd20576;
    data[ 3670] = -'sd19809;
    data[ 3671] =  'sd25178;
    data[ 3672] =  'sd12405;
    data[ 3673] = -'sd77006;
    data[ 3674] = -'sd47519;
    data[ 3675] = -'sd4951;
    data[ 3676] = -'sd34657;
    data[ 3677] = -'sd78758;
    data[ 3678] = -'sd59783;
    data[ 3679] =  'sd73042;
    data[ 3680] =  'sd19771;
    data[ 3681] = -'sd25444;
    data[ 3682] = -'sd14267;
    data[ 3683] =  'sd63972;
    data[ 3684] = -'sd43719;
    data[ 3685] =  'sd21649;
    data[ 3686] = -'sd12298;
    data[ 3687] =  'sd77755;
    data[ 3688] =  'sd52762;
    data[ 3689] =  'sd41652;
    data[ 3690] = -'sd36118;
    data[ 3691] =  'sd74856;
    data[ 3692] =  'sd32469;
    data[ 3693] =  'sd63442;
    data[ 3694] = -'sd47429;
    data[ 3695] = -'sd4321;
    data[ 3696] = -'sd30247;
    data[ 3697] = -'sd47888;
    data[ 3698] = -'sd7534;
    data[ 3699] = -'sd52738;
    data[ 3700] = -'sd41484;
    data[ 3701] =  'sd37294;
    data[ 3702] = -'sd66624;
    data[ 3703] =  'sd25155;
    data[ 3704] =  'sd12244;
    data[ 3705] = -'sd78133;
    data[ 3706] = -'sd55408;
    data[ 3707] = -'sd60174;
    data[ 3708] =  'sd70305;
    data[ 3709] =  'sd612;
    data[ 3710] =  'sd4284;
    data[ 3711] =  'sd29988;
    data[ 3712] =  'sd46075;
    data[ 3713] = -'sd5157;
    data[ 3714] = -'sd36099;
    data[ 3715] =  'sd74989;
    data[ 3716] =  'sd33400;
    data[ 3717] =  'sd69959;
    data[ 3718] = -'sd1810;
    data[ 3719] = -'sd12670;
    data[ 3720] =  'sd75151;
    data[ 3721] =  'sd34534;
    data[ 3722] =  'sd77897;
    data[ 3723] =  'sd53756;
    data[ 3724] =  'sd48610;
    data[ 3725] =  'sd12588;
    data[ 3726] = -'sd75725;
    data[ 3727] = -'sd38552;
    data[ 3728] =  'sd57818;
    data[ 3729] =  'sd77044;
    data[ 3730] =  'sd47785;
    data[ 3731] =  'sd6813;
    data[ 3732] =  'sd47691;
    data[ 3733] =  'sd6155;
    data[ 3734] =  'sd43085;
    data[ 3735] = -'sd26087;
    data[ 3736] = -'sd18768;
    data[ 3737] =  'sd32465;
    data[ 3738] =  'sd63414;
    data[ 3739] = -'sd47625;
    data[ 3740] = -'sd5693;
    data[ 3741] = -'sd39851;
    data[ 3742] =  'sd48725;
    data[ 3743] =  'sd13393;
    data[ 3744] = -'sd70090;
    data[ 3745] =  'sd893;
    data[ 3746] =  'sd6251;
    data[ 3747] =  'sd43757;
    data[ 3748] = -'sd21383;
    data[ 3749] =  'sd14160;
    data[ 3750] = -'sd64721;
    data[ 3751] =  'sd38476;
    data[ 3752] = -'sd58350;
    data[ 3753] = -'sd80768;
    data[ 3754] = -'sd73853;
    data[ 3755] = -'sd25448;
    data[ 3756] = -'sd14295;
    data[ 3757] =  'sd63776;
    data[ 3758] = -'sd45091;
    data[ 3759] =  'sd12045;
    data[ 3760] = -'sd79526;
    data[ 3761] = -'sd65159;
    data[ 3762] =  'sd35410;
    data[ 3763] = -'sd79812;
    data[ 3764] = -'sd67161;
    data[ 3765] =  'sd21396;
    data[ 3766] = -'sd14069;
    data[ 3767] =  'sd65358;
    data[ 3768] = -'sd34017;
    data[ 3769] = -'sd74278;
    data[ 3770] = -'sd28423;
    data[ 3771] = -'sd35120;
    data[ 3772] =  'sd81842;
    data[ 3773] =  'sd81371;
    data[ 3774] =  'sd78074;
    data[ 3775] =  'sd54995;
    data[ 3776] =  'sd57283;
    data[ 3777] =  'sd73299;
    data[ 3778] =  'sd21570;
    data[ 3779] = -'sd12851;
    data[ 3780] =  'sd73884;
    data[ 3781] =  'sd25665;
    data[ 3782] =  'sd15814;
    data[ 3783] = -'sd53143;
    data[ 3784] = -'sd44319;
    data[ 3785] =  'sd17449;
    data[ 3786] = -'sd41698;
    data[ 3787] =  'sd35796;
    data[ 3788] = -'sd77110;
    data[ 3789] = -'sd48247;
    data[ 3790] = -'sd10047;
    data[ 3791] = -'sd70329;
    data[ 3792] = -'sd780;
    data[ 3793] = -'sd5460;
    data[ 3794] = -'sd38220;
    data[ 3795] =  'sd60142;
    data[ 3796] = -'sd70529;
    data[ 3797] = -'sd2180;
    data[ 3798] = -'sd15260;
    data[ 3799] =  'sd57021;
    data[ 3800] =  'sd71465;
    data[ 3801] =  'sd8732;
    data[ 3802] =  'sd61124;
    data[ 3803] = -'sd63655;
    data[ 3804] =  'sd45938;
    data[ 3805] = -'sd6116;
    data[ 3806] = -'sd42812;
    data[ 3807] =  'sd27998;
    data[ 3808] =  'sd32145;
    data[ 3809] =  'sd61174;
    data[ 3810] = -'sd63305;
    data[ 3811] =  'sd48388;
    data[ 3812] =  'sd11034;
    data[ 3813] =  'sd77238;
    data[ 3814] =  'sd49143;
    data[ 3815] =  'sd16319;
    data[ 3816] = -'sd49608;
    data[ 3817] = -'sd19574;
    data[ 3818] =  'sd26823;
    data[ 3819] =  'sd23920;
    data[ 3820] =  'sd3599;
    data[ 3821] =  'sd25193;
    data[ 3822] =  'sd12510;
    data[ 3823] = -'sd76271;
    data[ 3824] = -'sd42374;
    data[ 3825] =  'sd31064;
    data[ 3826] =  'sd53607;
    data[ 3827] =  'sd47567;
    data[ 3828] =  'sd5287;
    data[ 3829] =  'sd37009;
    data[ 3830] = -'sd68619;
    data[ 3831] =  'sd11190;
    data[ 3832] =  'sd78330;
    data[ 3833] =  'sd56787;
    data[ 3834] =  'sd69827;
    data[ 3835] = -'sd2734;
    data[ 3836] = -'sd19138;
    data[ 3837] =  'sd29875;
    data[ 3838] =  'sd45284;
    data[ 3839] = -'sd10694;
    data[ 3840] = -'sd74858;
    data[ 3841] = -'sd32483;
    data[ 3842] = -'sd63540;
    data[ 3843] =  'sd46743;
    data[ 3844] = -'sd481;
    data[ 3845] = -'sd3367;
    data[ 3846] = -'sd23569;
    data[ 3847] = -'sd1142;
    data[ 3848] = -'sd7994;
    data[ 3849] = -'sd55958;
    data[ 3850] = -'sd64024;
    data[ 3851] =  'sd43355;
    data[ 3852] = -'sd24197;
    data[ 3853] = -'sd5538;
    data[ 3854] = -'sd38766;
    data[ 3855] =  'sd56320;
    data[ 3856] =  'sd66558;
    data[ 3857] = -'sd25617;
    data[ 3858] = -'sd15478;
    data[ 3859] =  'sd55495;
    data[ 3860] =  'sd60783;
    data[ 3861] = -'sd66042;
    data[ 3862] =  'sd29229;
    data[ 3863] =  'sd40762;
    data[ 3864] = -'sd42348;
    data[ 3865] =  'sd31246;
    data[ 3866] =  'sd54881;
    data[ 3867] =  'sd56485;
    data[ 3868] =  'sd67713;
    data[ 3869] = -'sd17532;
    data[ 3870] =  'sd41117;
    data[ 3871] = -'sd39863;
    data[ 3872] =  'sd48641;
    data[ 3873] =  'sd12805;
    data[ 3874] = -'sd74206;
    data[ 3875] = -'sd27919;
    data[ 3876] = -'sd31592;
    data[ 3877] = -'sd57303;
    data[ 3878] = -'sd73439;
    data[ 3879] = -'sd22550;
    data[ 3880] =  'sd5991;
    data[ 3881] =  'sd41937;
    data[ 3882] = -'sd34123;
    data[ 3883] = -'sd75020;
    data[ 3884] = -'sd33617;
    data[ 3885] = -'sd71478;
    data[ 3886] = -'sd8823;
    data[ 3887] = -'sd61761;
    data[ 3888] =  'sd59196;
    data[ 3889] = -'sd77151;
    data[ 3890] = -'sd48534;
    data[ 3891] = -'sd12056;
    data[ 3892] =  'sd79449;
    data[ 3893] =  'sd64620;
    data[ 3894] = -'sd39183;
    data[ 3895] =  'sd53401;
    data[ 3896] =  'sd46125;
    data[ 3897] = -'sd4807;
    data[ 3898] = -'sd33649;
    data[ 3899] = -'sd71702;
    data[ 3900] = -'sd10391;
    data[ 3901] = -'sd72737;
    data[ 3902] = -'sd17636;
    data[ 3903] =  'sd40389;
    data[ 3904] = -'sd44959;
    data[ 3905] =  'sd12969;
    data[ 3906] = -'sd73058;
    data[ 3907] = -'sd19883;
    data[ 3908] =  'sd24660;
    data[ 3909] =  'sd8779;
    data[ 3910] =  'sd61453;
    data[ 3911] = -'sd61352;
    data[ 3912] =  'sd62059;
    data[ 3913] = -'sd57110;
    data[ 3914] = -'sd72088;
    data[ 3915] = -'sd13093;
    data[ 3916] =  'sd72190;
    data[ 3917] =  'sd13807;
    data[ 3918] = -'sd67192;
    data[ 3919] =  'sd21179;
    data[ 3920] = -'sd15588;
    data[ 3921] =  'sd54725;
    data[ 3922] =  'sd55393;
    data[ 3923] =  'sd60069;
    data[ 3924] = -'sd71040;
    data[ 3925] = -'sd5757;
    data[ 3926] = -'sd40299;
    data[ 3927] =  'sd45589;
    data[ 3928] = -'sd8559;
    data[ 3929] = -'sd59913;
    data[ 3930] =  'sd72132;
    data[ 3931] =  'sd13401;
    data[ 3932] = -'sd70034;
    data[ 3933] =  'sd1285;
    data[ 3934] =  'sd8995;
    data[ 3935] =  'sd62965;
    data[ 3936] = -'sd50768;
    data[ 3937] = -'sd27694;
    data[ 3938] = -'sd30017;
    data[ 3939] = -'sd46278;
    data[ 3940] =  'sd3736;
    data[ 3941] =  'sd26152;
    data[ 3942] =  'sd19223;
    data[ 3943] = -'sd29280;
    data[ 3944] = -'sd41119;
    data[ 3945] =  'sd39849;
    data[ 3946] = -'sd48739;
    data[ 3947] = -'sd13491;
    data[ 3948] =  'sd69404;
    data[ 3949] = -'sd5695;
    data[ 3950] = -'sd39865;
    data[ 3951] =  'sd48627;
    data[ 3952] =  'sd12707;
    data[ 3953] = -'sd74892;
    data[ 3954] = -'sd32721;
    data[ 3955] = -'sd65206;
    data[ 3956] =  'sd35081;
    data[ 3957] =  'sd81726;
    data[ 3958] =  'sd80559;
    data[ 3959] =  'sd72390;
    data[ 3960] =  'sd15207;
    data[ 3961] = -'sd57392;
    data[ 3962] = -'sd74062;
    data[ 3963] = -'sd26911;
    data[ 3964] = -'sd24536;
    data[ 3965] = -'sd7911;
    data[ 3966] = -'sd55377;
    data[ 3967] = -'sd59957;
    data[ 3968] =  'sd71824;
    data[ 3969] =  'sd11245;
    data[ 3970] =  'sd78715;
    data[ 3971] =  'sd59482;
    data[ 3972] = -'sd75149;
    data[ 3973] = -'sd34520;
    data[ 3974] = -'sd77799;
    data[ 3975] = -'sd53070;
    data[ 3976] = -'sd43808;
    data[ 3977] =  'sd21026;
    data[ 3978] = -'sd16659;
    data[ 3979] =  'sd47228;
    data[ 3980] =  'sd2914;
    data[ 3981] =  'sd20398;
    data[ 3982] = -'sd21055;
    data[ 3983] =  'sd16456;
    data[ 3984] = -'sd48649;
    data[ 3985] = -'sd12861;
    data[ 3986] =  'sd73814;
    data[ 3987] =  'sd25175;
    data[ 3988] =  'sd12384;
    data[ 3989] = -'sd77153;
    data[ 3990] = -'sd48548;
    data[ 3991] = -'sd12154;
    data[ 3992] =  'sd78763;
    data[ 3993] =  'sd59818;
    data[ 3994] = -'sd72797;
    data[ 3995] = -'sd18056;
    data[ 3996] =  'sd37449;
    data[ 3997] = -'sd65539;
    data[ 3998] =  'sd32750;
    data[ 3999] =  'sd65409;
    data[ 4000] = -'sd33660;
    data[ 4001] = -'sd71779;
    data[ 4002] = -'sd10930;
    data[ 4003] = -'sd76510;
    data[ 4004] = -'sd44047;
    data[ 4005] =  'sd19353;
    data[ 4006] = -'sd28370;
    data[ 4007] = -'sd34749;
    data[ 4008] = -'sd79402;
    data[ 4009] = -'sd64291;
    data[ 4010] =  'sd41486;
    data[ 4011] = -'sd37280;
    data[ 4012] =  'sd66722;
    data[ 4013] = -'sd24469;
    data[ 4014] = -'sd7442;
    data[ 4015] = -'sd52094;
    data[ 4016] = -'sd36976;
    data[ 4017] =  'sd68850;
    data[ 4018] = -'sd9573;
    data[ 4019] = -'sd67011;
    data[ 4020] =  'sd22446;
    data[ 4021] = -'sd6719;
    data[ 4022] = -'sd47033;
    data[ 4023] = -'sd1549;
    data[ 4024] = -'sd10843;
    data[ 4025] = -'sd75901;
    data[ 4026] = -'sd39784;
    data[ 4027] =  'sd49194;
    data[ 4028] =  'sd16676;
    data[ 4029] = -'sd47109;
    data[ 4030] = -'sd2081;
    data[ 4031] = -'sd14567;
    data[ 4032] =  'sd61872;
    data[ 4033] = -'sd58419;
    data[ 4034] = -'sd81251;
    data[ 4035] = -'sd77234;
    data[ 4036] = -'sd49115;
    data[ 4037] = -'sd16123;
    data[ 4038] =  'sd50980;
    data[ 4039] =  'sd29178;
    data[ 4040] =  'sd40405;
    data[ 4041] = -'sd44847;
    data[ 4042] =  'sd13753;
    data[ 4043] = -'sd67570;
    data[ 4044] =  'sd18533;
    data[ 4045] = -'sd34110;
    data[ 4046] = -'sd74929;
    data[ 4047] = -'sd32980;
    data[ 4048] = -'sd67019;
    data[ 4049] =  'sd22390;
    data[ 4050] = -'sd7111;
    data[ 4051] = -'sd49777;
    data[ 4052] = -'sd20757;
    data[ 4053] =  'sd18542;
    data[ 4054] = -'sd34047;
    data[ 4055] = -'sd74488;
    data[ 4056] = -'sd29893;
    data[ 4057] = -'sd45410;
    data[ 4058] =  'sd9812;
    data[ 4059] =  'sd68684;
    data[ 4060] = -'sd10735;
    data[ 4061] = -'sd75145;
    data[ 4062] = -'sd34492;
    data[ 4063] = -'sd77603;
    data[ 4064] = -'sd51698;
    data[ 4065] = -'sd34204;
    data[ 4066] = -'sd75587;
    data[ 4067] = -'sd37586;
    data[ 4068] =  'sd64580;
    data[ 4069] = -'sd39463;
    data[ 4070] =  'sd51441;
    data[ 4071] =  'sd32405;
    data[ 4072] =  'sd62994;
    data[ 4073] = -'sd50565;
    data[ 4074] = -'sd26273;
    data[ 4075] = -'sd20070;
    data[ 4076] =  'sd23351;
    data[ 4077] = -'sd384;
    data[ 4078] = -'sd2688;
    data[ 4079] = -'sd18816;
    data[ 4080] =  'sd32129;
    data[ 4081] =  'sd61062;
    data[ 4082] = -'sd64089;
    data[ 4083] =  'sd42900;
    data[ 4084] = -'sd27382;
    data[ 4085] = -'sd27833;
    data[ 4086] = -'sd30990;
    data[ 4087] = -'sd53089;
    data[ 4088] = -'sd43941;
    data[ 4089] =  'sd20095;
    data[ 4090] = -'sd23176;
    data[ 4091] =  'sd1609;
    data[ 4092] =  'sd11263;
    data[ 4093] =  'sd78841;
    data[ 4094] =  'sd60364;
    data[ 4095] = -'sd68975;
    data[ 4096] =  'sd8698;
    data[ 4097] =  'sd60886;
    data[ 4098] = -'sd65321;
    data[ 4099] =  'sd34276;
    data[ 4100] =  'sd76091;
    data[ 4101] =  'sd41114;
    data[ 4102] = -'sd39884;
    data[ 4103] =  'sd48494;
    data[ 4104] =  'sd11776;
    data[ 4105] = -'sd81409;
    data[ 4106] = -'sd78340;
    data[ 4107] = -'sd56857;
    data[ 4108] = -'sd70317;
    data[ 4109] = -'sd696;
    data[ 4110] = -'sd4872;
    data[ 4111] = -'sd34104;
    data[ 4112] = -'sd74887;
    data[ 4113] = -'sd32686;
    data[ 4114] = -'sd64961;
    data[ 4115] =  'sd36796;
    data[ 4116] = -'sd70110;
    data[ 4117] =  'sd753;
    data[ 4118] =  'sd5271;
    data[ 4119] =  'sd36897;
    data[ 4120] = -'sd69403;
    data[ 4121] =  'sd5702;
    data[ 4122] =  'sd39914;
    data[ 4123] = -'sd48284;
    data[ 4124] = -'sd10306;
    data[ 4125] = -'sd72142;
    data[ 4126] = -'sd13471;
    data[ 4127] =  'sd69544;
    data[ 4128] = -'sd4715;
    data[ 4129] = -'sd33005;
    data[ 4130] = -'sd67194;
    data[ 4131] =  'sd21165;
    data[ 4132] = -'sd15686;
    data[ 4133] =  'sd54039;
    data[ 4134] =  'sd50591;
    data[ 4135] =  'sd26455;
    data[ 4136] =  'sd21344;
    data[ 4137] = -'sd14433;
    data[ 4138] =  'sd62810;
    data[ 4139] = -'sd51853;
    data[ 4140] = -'sd35289;
    data[ 4141] =  'sd80659;
    data[ 4142] =  'sd73090;
    data[ 4143] =  'sd20107;
    data[ 4144] = -'sd23092;
    data[ 4145] =  'sd2197;
    data[ 4146] =  'sd15379;
    data[ 4147] = -'sd56188;
    data[ 4148] = -'sd65634;
    data[ 4149] =  'sd32085;
    data[ 4150] =  'sd60754;
    data[ 4151] = -'sd66245;
    data[ 4152] =  'sd27808;
    data[ 4153] =  'sd30815;
    data[ 4154] =  'sd51864;
    data[ 4155] =  'sd35366;
    data[ 4156] = -'sd80120;
    data[ 4157] = -'sd69317;
    data[ 4158] =  'sd6304;
    data[ 4159] =  'sd44128;
    data[ 4160] = -'sd18786;
    data[ 4161] =  'sd32339;
    data[ 4162] =  'sd62532;
    data[ 4163] = -'sd53799;
    data[ 4164] = -'sd48911;
    data[ 4165] = -'sd14695;
    data[ 4166] =  'sd60976;
    data[ 4167] = -'sd64691;
    data[ 4168] =  'sd38686;
    data[ 4169] = -'sd56880;
    data[ 4170] = -'sd70478;
    data[ 4171] = -'sd1823;
    data[ 4172] = -'sd12761;
    data[ 4173] =  'sd74514;
    data[ 4174] =  'sd30075;
    data[ 4175] =  'sd46684;
    data[ 4176] = -'sd894;
    data[ 4177] = -'sd6258;
    data[ 4178] = -'sd43806;
    data[ 4179] =  'sd21040;
    data[ 4180] = -'sd16561;
    data[ 4181] =  'sd47914;
    data[ 4182] =  'sd7716;
    data[ 4183] =  'sd54012;
    data[ 4184] =  'sd50402;
    data[ 4185] =  'sd25132;
    data[ 4186] =  'sd12083;
    data[ 4187] = -'sd79260;
    data[ 4188] = -'sd63297;
    data[ 4189] =  'sd48444;
    data[ 4190] =  'sd11426;
    data[ 4191] =  'sd79982;
    data[ 4192] =  'sd68351;
    data[ 4193] = -'sd13066;
    data[ 4194] =  'sd72379;
    data[ 4195] =  'sd15130;
    data[ 4196] = -'sd57931;
    data[ 4197] = -'sd77835;
    data[ 4198] = -'sd53322;
    data[ 4199] = -'sd45572;
    data[ 4200] =  'sd8678;
    data[ 4201] =  'sd60746;
    data[ 4202] = -'sd66301;
    data[ 4203] =  'sd27416;
    data[ 4204] =  'sd28071;
    data[ 4205] =  'sd32656;
    data[ 4206] =  'sd64751;
    data[ 4207] = -'sd38266;
    data[ 4208] =  'sd59820;
    data[ 4209] = -'sd72783;
    data[ 4210] = -'sd17958;
    data[ 4211] =  'sd38135;
    data[ 4212] = -'sd60737;
    data[ 4213] =  'sd66364;
    data[ 4214] = -'sd26975;
    data[ 4215] = -'sd24984;
    data[ 4216] = -'sd11047;
    data[ 4217] = -'sd77329;
    data[ 4218] = -'sd49780;
    data[ 4219] = -'sd20778;
    data[ 4220] =  'sd18395;
    data[ 4221] = -'sd35076;
    data[ 4222] = -'sd81691;
    data[ 4223] = -'sd80314;
    data[ 4224] = -'sd70675;
    data[ 4225] = -'sd3202;
    data[ 4226] = -'sd22414;
    data[ 4227] =  'sd6943;
    data[ 4228] =  'sd48601;
    data[ 4229] =  'sd12525;
    data[ 4230] = -'sd76166;
    data[ 4231] = -'sd41639;
    data[ 4232] =  'sd36209;
    data[ 4233] = -'sd74219;
    data[ 4234] = -'sd28010;
    data[ 4235] = -'sd32229;
    data[ 4236] = -'sd61762;
    data[ 4237] =  'sd59189;
    data[ 4238] = -'sd77200;
    data[ 4239] = -'sd48877;
    data[ 4240] = -'sd14457;
    data[ 4241] =  'sd62642;
    data[ 4242] = -'sd53029;
    data[ 4243] = -'sd43521;
    data[ 4244] =  'sd23035;
    data[ 4245] = -'sd2596;
    data[ 4246] = -'sd18172;
    data[ 4247] =  'sd36637;
    data[ 4248] = -'sd71223;
    data[ 4249] = -'sd7038;
    data[ 4250] = -'sd49266;
    data[ 4251] = -'sd17180;
    data[ 4252] =  'sd43581;
    data[ 4253] = -'sd22615;
    data[ 4254] =  'sd5536;
    data[ 4255] =  'sd38752;
    data[ 4256] = -'sd56418;
    data[ 4257] = -'sd67244;
    data[ 4258] =  'sd20815;
    data[ 4259] = -'sd18136;
    data[ 4260] =  'sd36889;
    data[ 4261] = -'sd69459;
    data[ 4262] =  'sd5310;
    data[ 4263] =  'sd37170;
    data[ 4264] = -'sd67492;
    data[ 4265] =  'sd19079;
    data[ 4266] = -'sd30288;
    data[ 4267] = -'sd48175;
    data[ 4268] = -'sd9543;
    data[ 4269] = -'sd66801;
    data[ 4270] =  'sd23916;
    data[ 4271] =  'sd3571;
    data[ 4272] =  'sd24997;
    data[ 4273] =  'sd11138;
    data[ 4274] =  'sd77966;
    data[ 4275] =  'sd54239;
    data[ 4276] =  'sd51991;
    data[ 4277] =  'sd36255;
    data[ 4278] = -'sd73897;
    data[ 4279] = -'sd25756;
    data[ 4280] = -'sd16451;
    data[ 4281] =  'sd48684;
    data[ 4282] =  'sd13106;
    data[ 4283] = -'sd72099;
    data[ 4284] = -'sd13170;
    data[ 4285] =  'sd71651;
    data[ 4286] =  'sd10034;
    data[ 4287] =  'sd70238;
    data[ 4288] =  'sd143;
    data[ 4289] =  'sd1001;
    data[ 4290] =  'sd7007;
    data[ 4291] =  'sd49049;
    data[ 4292] =  'sd15661;
    data[ 4293] = -'sd54214;
    data[ 4294] = -'sd51816;
    data[ 4295] = -'sd35030;
    data[ 4296] = -'sd81369;
    data[ 4297] = -'sd78060;
    data[ 4298] = -'sd54897;
    data[ 4299] = -'sd56597;
    data[ 4300] = -'sd68497;
    data[ 4301] =  'sd12044;
    data[ 4302] = -'sd79533;
    data[ 4303] = -'sd65208;
    data[ 4304] =  'sd35067;
    data[ 4305] =  'sd81628;
    data[ 4306] =  'sd79873;
    data[ 4307] =  'sd67588;
    data[ 4308] = -'sd18407;
    data[ 4309] =  'sd34992;
    data[ 4310] =  'sd81103;
    data[ 4311] =  'sd76198;
    data[ 4312] =  'sd41863;
    data[ 4313] = -'sd34641;
    data[ 4314] = -'sd78646;
    data[ 4315] = -'sd58999;
    data[ 4316] =  'sd78530;
    data[ 4317] =  'sd58187;
    data[ 4318] =  'sd79627;
    data[ 4319] =  'sd65866;
    data[ 4320] = -'sd30461;
    data[ 4321] = -'sd49386;
    data[ 4322] = -'sd18020;
    data[ 4323] =  'sd37701;
    data[ 4324] = -'sd63775;
    data[ 4325] =  'sd45098;
    data[ 4326] = -'sd11996;
    data[ 4327] =  'sd79869;
    data[ 4328] =  'sd67560;
    data[ 4329] = -'sd18603;
    data[ 4330] =  'sd33620;
    data[ 4331] =  'sd71499;
    data[ 4332] =  'sd8970;
    data[ 4333] =  'sd62790;
    data[ 4334] = -'sd51993;
    data[ 4335] = -'sd36269;
    data[ 4336] =  'sd73799;
    data[ 4337] =  'sd25070;
    data[ 4338] =  'sd11649;
    data[ 4339] =  'sd81543;
    data[ 4340] =  'sd79278;
    data[ 4341] =  'sd63423;
    data[ 4342] = -'sd47562;
    data[ 4343] = -'sd5252;
    data[ 4344] = -'sd36764;
    data[ 4345] =  'sd70334;
    data[ 4346] =  'sd815;
    data[ 4347] =  'sd5705;
    data[ 4348] =  'sd39935;
    data[ 4349] = -'sd48137;
    data[ 4350] = -'sd9277;
    data[ 4351] = -'sd64939;
    data[ 4352] =  'sd36950;
    data[ 4353] = -'sd69032;
    data[ 4354] =  'sd8299;
    data[ 4355] =  'sd58093;
    data[ 4356] =  'sd78969;
    data[ 4357] =  'sd61260;
    data[ 4358] = -'sd62703;
    data[ 4359] =  'sd52602;
    data[ 4360] =  'sd40532;
    data[ 4361] = -'sd43958;
    data[ 4362] =  'sd19976;
    data[ 4363] = -'sd24009;
    data[ 4364] = -'sd4222;
    data[ 4365] = -'sd29554;
    data[ 4366] = -'sd43037;
    data[ 4367] =  'sd26423;
    data[ 4368] =  'sd21120;
    data[ 4369] = -'sd16001;
    data[ 4370] =  'sd51834;
    data[ 4371] =  'sd35156;
    data[ 4372] = -'sd81590;
    data[ 4373] = -'sd79607;
    data[ 4374] = -'sd65726;
    data[ 4375] =  'sd31441;
    data[ 4376] =  'sd56246;
    data[ 4377] =  'sd66040;
    data[ 4378] = -'sd29243;
    data[ 4379] = -'sd40860;
    data[ 4380] =  'sd41662;
    data[ 4381] = -'sd36048;
    data[ 4382] =  'sd75346;
    data[ 4383] =  'sd35899;
    data[ 4384] = -'sd76389;
    data[ 4385] = -'sd43200;
    data[ 4386] =  'sd25282;
    data[ 4387] =  'sd13133;
    data[ 4388] = -'sd71910;
    data[ 4389] = -'sd11847;
    data[ 4390] =  'sd80912;
    data[ 4391] =  'sd74861;
    data[ 4392] =  'sd32504;
    data[ 4393] =  'sd63687;
    data[ 4394] = -'sd45714;
    data[ 4395] =  'sd7684;
    data[ 4396] =  'sd53788;
    data[ 4397] =  'sd48834;
    data[ 4398] =  'sd14156;
    data[ 4399] = -'sd64749;
    data[ 4400] =  'sd38280;
    data[ 4401] = -'sd59722;
    data[ 4402] =  'sd73469;
    data[ 4403] =  'sd22760;
    data[ 4404] = -'sd4521;
    data[ 4405] = -'sd31647;
    data[ 4406] = -'sd57688;
    data[ 4407] = -'sd76134;
    data[ 4408] = -'sd41415;
    data[ 4409] =  'sd37777;
    data[ 4410] = -'sd63243;
    data[ 4411] =  'sd48822;
    data[ 4412] =  'sd14072;
    data[ 4413] = -'sd65337;
    data[ 4414] =  'sd34164;
    data[ 4415] =  'sd75307;
    data[ 4416] =  'sd35626;
    data[ 4417] = -'sd78300;
    data[ 4418] = -'sd56577;
    data[ 4419] = -'sd68357;
    data[ 4420] =  'sd13024;
    data[ 4421] = -'sd72673;
    data[ 4422] = -'sd17188;
    data[ 4423] =  'sd43525;
    data[ 4424] = -'sd23007;
    data[ 4425] =  'sd2792;
    data[ 4426] =  'sd19544;
    data[ 4427] = -'sd27033;
    data[ 4428] = -'sd25390;
    data[ 4429] = -'sd13889;
    data[ 4430] =  'sd66618;
    data[ 4431] = -'sd25197;
    data[ 4432] = -'sd12538;
    data[ 4433] =  'sd76075;
    data[ 4434] =  'sd41002;
    data[ 4435] = -'sd40668;
    data[ 4436] =  'sd43006;
    data[ 4437] = -'sd26640;
    data[ 4438] = -'sd22639;
    data[ 4439] =  'sd5368;
    data[ 4440] =  'sd37576;
    data[ 4441] = -'sd64650;
    data[ 4442] =  'sd38973;
    data[ 4443] = -'sd54871;
    data[ 4444] = -'sd56415;
    data[ 4445] = -'sd67223;
    data[ 4446] =  'sd20962;
    data[ 4447] = -'sd17107;
    data[ 4448] =  'sd44092;
    data[ 4449] = -'sd19038;
    data[ 4450] =  'sd30575;
    data[ 4451] =  'sd50184;
    data[ 4452] =  'sd23606;
    data[ 4453] =  'sd1401;
    data[ 4454] =  'sd9807;
    data[ 4455] =  'sd68649;
    data[ 4456] = -'sd10980;
    data[ 4457] = -'sd76860;
    data[ 4458] = -'sd46497;
    data[ 4459] =  'sd2203;
    data[ 4460] =  'sd15421;
    data[ 4461] = -'sd55894;
    data[ 4462] = -'sd63576;
    data[ 4463] =  'sd46491;
    data[ 4464] = -'sd2245;
    data[ 4465] = -'sd15715;
    data[ 4466] =  'sd53836;
    data[ 4467] =  'sd49170;
    data[ 4468] =  'sd16508;
    data[ 4469] = -'sd48285;
    data[ 4470] = -'sd10313;
    data[ 4471] = -'sd72191;
    data[ 4472] = -'sd13814;
    data[ 4473] =  'sd67143;
    data[ 4474] = -'sd21522;
    data[ 4475] =  'sd13187;
    data[ 4476] = -'sd71532;
    data[ 4477] = -'sd9201;
    data[ 4478] = -'sd64407;
    data[ 4479] =  'sd40674;
    data[ 4480] = -'sd42964;
    data[ 4481] =  'sd26934;
    data[ 4482] =  'sd24697;
    data[ 4483] =  'sd9038;
    data[ 4484] =  'sd63266;
    data[ 4485] = -'sd48661;
    data[ 4486] = -'sd12945;
    data[ 4487] =  'sd73226;
    data[ 4488] =  'sd21059;
    data[ 4489] = -'sd16428;
    data[ 4490] =  'sd48845;
    data[ 4491] =  'sd14233;
    data[ 4492] = -'sd64210;
    data[ 4493] =  'sd42053;
    data[ 4494] = -'sd33311;
    data[ 4495] = -'sd69336;
    data[ 4496] =  'sd6171;
    data[ 4497] =  'sd43197;
    data[ 4498] = -'sd25303;
    data[ 4499] = -'sd13280;
    data[ 4500] =  'sd70881;
    data[ 4501] =  'sd4644;
    data[ 4502] =  'sd32508;
    data[ 4503] =  'sd63715;
    data[ 4504] = -'sd45518;
    data[ 4505] =  'sd9056;
    data[ 4506] =  'sd63392;
    data[ 4507] = -'sd47779;
    data[ 4508] = -'sd6771;
    data[ 4509] = -'sd47397;
    data[ 4510] = -'sd4097;
    data[ 4511] = -'sd28679;
    data[ 4512] = -'sd36912;
    data[ 4513] =  'sd69298;
    data[ 4514] = -'sd6437;
    data[ 4515] = -'sd45059;
    data[ 4516] =  'sd12269;
    data[ 4517] = -'sd77958;
    data[ 4518] = -'sd54183;
    data[ 4519] = -'sd51599;
    data[ 4520] = -'sd33511;
    data[ 4521] = -'sd70736;
    data[ 4522] = -'sd3629;
    data[ 4523] = -'sd25403;
    data[ 4524] = -'sd13980;
    data[ 4525] =  'sd65981;
    data[ 4526] = -'sd29656;
    data[ 4527] = -'sd43751;
    data[ 4528] =  'sd21425;
    data[ 4529] = -'sd13866;
    data[ 4530] =  'sd66779;
    data[ 4531] = -'sd24070;
    data[ 4532] = -'sd4649;
    data[ 4533] = -'sd32543;
    data[ 4534] = -'sd63960;
    data[ 4535] =  'sd43803;
    data[ 4536] = -'sd21061;
    data[ 4537] =  'sd16414;
    data[ 4538] = -'sd48943;
    data[ 4539] = -'sd14919;
    data[ 4540] =  'sd59408;
    data[ 4541] = -'sd75667;
    data[ 4542] = -'sd38146;
    data[ 4543] =  'sd60660;
    data[ 4544] = -'sd66903;
    data[ 4545] =  'sd23202;
    data[ 4546] = -'sd1427;
    data[ 4547] = -'sd9989;
    data[ 4548] = -'sd69923;
    data[ 4549] =  'sd2062;
    data[ 4550] =  'sd14434;
    data[ 4551] = -'sd62803;
    data[ 4552] =  'sd51902;
    data[ 4553] =  'sd35632;
    data[ 4554] = -'sd78258;
    data[ 4555] = -'sd56283;
    data[ 4556] = -'sd66299;
    data[ 4557] =  'sd27430;
    data[ 4558] =  'sd28169;
    data[ 4559] =  'sd33342;
    data[ 4560] =  'sd69553;
    data[ 4561] = -'sd4652;
    data[ 4562] = -'sd32564;
    data[ 4563] = -'sd64107;
    data[ 4564] =  'sd42774;
    data[ 4565] = -'sd28264;
    data[ 4566] = -'sd34007;
    data[ 4567] = -'sd74208;
    data[ 4568] = -'sd27933;
    data[ 4569] = -'sd31690;
    data[ 4570] = -'sd57989;
    data[ 4571] = -'sd78241;
    data[ 4572] = -'sd56164;
    data[ 4573] = -'sd65466;
    data[ 4574] =  'sd33261;
    data[ 4575] =  'sd68986;
    data[ 4576] = -'sd8621;
    data[ 4577] = -'sd60347;
    data[ 4578] =  'sd69094;
    data[ 4579] = -'sd7865;
    data[ 4580] = -'sd55055;
    data[ 4581] = -'sd57703;
    data[ 4582] = -'sd76239;
    data[ 4583] = -'sd42150;
    data[ 4584] =  'sd32632;
    data[ 4585] =  'sd64583;
    data[ 4586] = -'sd39442;
    data[ 4587] =  'sd51588;
    data[ 4588] =  'sd33434;
    data[ 4589] =  'sd70197;
    data[ 4590] = -'sd144;
    data[ 4591] = -'sd1008;
    data[ 4592] = -'sd7056;
    data[ 4593] = -'sd49392;
    data[ 4594] = -'sd18062;
    data[ 4595] =  'sd37407;
    data[ 4596] = -'sd65833;
    data[ 4597] =  'sd30692;
    data[ 4598] =  'sd51003;
    data[ 4599] =  'sd29339;
    data[ 4600] =  'sd41532;
    data[ 4601] = -'sd36958;
    data[ 4602] =  'sd68976;
    data[ 4603] = -'sd8691;
    data[ 4604] = -'sd60837;
    data[ 4605] =  'sd65664;
    data[ 4606] = -'sd31875;
    data[ 4607] = -'sd59284;
    data[ 4608] =  'sd76535;
    data[ 4609] =  'sd44222;
    data[ 4610] = -'sd18128;
    data[ 4611] =  'sd36945;
    data[ 4612] = -'sd69067;
    data[ 4613] =  'sd8054;
    data[ 4614] =  'sd56378;
    data[ 4615] =  'sd66964;
    data[ 4616] = -'sd22775;
    data[ 4617] =  'sd4416;
    data[ 4618] =  'sd30912;
    data[ 4619] =  'sd52543;
    data[ 4620] =  'sd40119;
    data[ 4621] = -'sd46849;
    data[ 4622] = -'sd261;
    data[ 4623] = -'sd1827;
    data[ 4624] = -'sd12789;
    data[ 4625] =  'sd74318;
    data[ 4626] =  'sd28703;
    data[ 4627] =  'sd37080;
    data[ 4628] = -'sd68122;
    data[ 4629] =  'sd14669;
    data[ 4630] = -'sd61158;
    data[ 4631] =  'sd63417;
    data[ 4632] = -'sd47604;
    data[ 4633] = -'sd5546;
    data[ 4634] = -'sd38822;
    data[ 4635] =  'sd55928;
    data[ 4636] =  'sd63814;
    data[ 4637] = -'sd44825;
    data[ 4638] =  'sd13907;
    data[ 4639] = -'sd66492;
    data[ 4640] =  'sd26079;
    data[ 4641] =  'sd18712;
    data[ 4642] = -'sd32857;
    data[ 4643] = -'sd66158;
    data[ 4644] =  'sd28417;
    data[ 4645] =  'sd35078;
    data[ 4646] =  'sd81705;
    data[ 4647] =  'sd80412;
    data[ 4648] =  'sd71361;
    data[ 4649] =  'sd8004;
    data[ 4650] =  'sd56028;
    data[ 4651] =  'sd64514;
    data[ 4652] = -'sd39925;
    data[ 4653] =  'sd48207;
    data[ 4654] =  'sd9767;
    data[ 4655] =  'sd68369;
    data[ 4656] = -'sd12940;
    data[ 4657] =  'sd73261;
    data[ 4658] =  'sd21304;
    data[ 4659] = -'sd14713;
    data[ 4660] =  'sd60850;
    data[ 4661] = -'sd65573;
    data[ 4662] =  'sd32512;
    data[ 4663] =  'sd63743;
    data[ 4664] = -'sd45322;
    data[ 4665] =  'sd10428;
    data[ 4666] =  'sd72996;
    data[ 4667] =  'sd19449;
    data[ 4668] = -'sd27698;
    data[ 4669] = -'sd30045;
    data[ 4670] = -'sd46474;
    data[ 4671] =  'sd2364;
    data[ 4672] =  'sd16548;
    data[ 4673] = -'sd48005;
    data[ 4674] = -'sd8353;
    data[ 4675] = -'sd58471;
    data[ 4676] = -'sd81615;
    data[ 4677] = -'sd79782;
    data[ 4678] = -'sd66951;
    data[ 4679] =  'sd22866;
    data[ 4680] = -'sd3779;
    data[ 4681] = -'sd26453;
    data[ 4682] = -'sd21330;
    data[ 4683] =  'sd14531;
    data[ 4684] = -'sd62124;
    data[ 4685] =  'sd56655;
    data[ 4686] =  'sd68903;
    data[ 4687] = -'sd9202;
    data[ 4688] = -'sd64414;
    data[ 4689] =  'sd40625;
    data[ 4690] = -'sd43307;
    data[ 4691] =  'sd24533;
    data[ 4692] =  'sd7890;
    data[ 4693] =  'sd55230;
    data[ 4694] =  'sd58928;
    data[ 4695] = -'sd79027;
    data[ 4696] = -'sd61666;
    data[ 4697] =  'sd59861;
    data[ 4698] = -'sd72496;
    data[ 4699] = -'sd15949;
    data[ 4700] =  'sd52198;
    data[ 4701] =  'sd37704;
    data[ 4702] = -'sd63754;
    data[ 4703] =  'sd45245;
    data[ 4704] = -'sd10967;
    data[ 4705] = -'sd76769;
    data[ 4706] = -'sd45860;
    data[ 4707] =  'sd6662;
    data[ 4708] =  'sd46634;
    data[ 4709] = -'sd1244;
    data[ 4710] = -'sd8708;
    data[ 4711] = -'sd60956;
    data[ 4712] =  'sd64831;
    data[ 4713] = -'sd37706;
    data[ 4714] =  'sd63740;
    data[ 4715] = -'sd45343;
    data[ 4716] =  'sd10281;
    data[ 4717] =  'sd71967;
    data[ 4718] =  'sd12246;
    data[ 4719] = -'sd78119;
    data[ 4720] = -'sd55310;
    data[ 4721] = -'sd59488;
    data[ 4722] =  'sd75107;
    data[ 4723] =  'sd34226;
    data[ 4724] =  'sd75741;
    data[ 4725] =  'sd38664;
    data[ 4726] = -'sd57034;
    data[ 4727] = -'sd71556;
    data[ 4728] = -'sd9369;
    data[ 4729] = -'sd65583;
    data[ 4730] =  'sd32442;
    data[ 4731] =  'sd63253;
    data[ 4732] = -'sd48752;
    data[ 4733] = -'sd13582;
    data[ 4734] =  'sd68767;
    data[ 4735] = -'sd10154;
    data[ 4736] = -'sd71078;
    data[ 4737] = -'sd6023;
    data[ 4738] = -'sd42161;
    data[ 4739] =  'sd32555;
    data[ 4740] =  'sd64044;
    data[ 4741] = -'sd43215;
    data[ 4742] =  'sd25177;
    data[ 4743] =  'sd12398;
    data[ 4744] = -'sd77055;
    data[ 4745] = -'sd47862;
    data[ 4746] = -'sd7352;
    data[ 4747] = -'sd51464;
    data[ 4748] = -'sd32566;
    data[ 4749] = -'sd64121;
    data[ 4750] =  'sd42676;
    data[ 4751] = -'sd28950;
    data[ 4752] = -'sd38809;
    data[ 4753] =  'sd56019;
    data[ 4754] =  'sd64451;
    data[ 4755] = -'sd40366;
    data[ 4756] =  'sd45120;
    data[ 4757] = -'sd11842;
    data[ 4758] =  'sd80947;
    data[ 4759] =  'sd75106;
    data[ 4760] =  'sd34219;
    data[ 4761] =  'sd75692;
    data[ 4762] =  'sd38321;
    data[ 4763] = -'sd59435;
    data[ 4764] =  'sd75478;
    data[ 4765] =  'sd36823;
    data[ 4766] = -'sd69921;
    data[ 4767] =  'sd2076;
    data[ 4768] =  'sd14532;
    data[ 4769] = -'sd62117;
    data[ 4770] =  'sd56704;
    data[ 4771] =  'sd69246;
    data[ 4772] = -'sd6801;
    data[ 4773] = -'sd47607;
    data[ 4774] = -'sd5567;
    data[ 4775] = -'sd38969;
    data[ 4776] =  'sd54899;
    data[ 4777] =  'sd56611;
    data[ 4778] =  'sd68595;
    data[ 4779] = -'sd11358;
    data[ 4780] = -'sd79506;
    data[ 4781] = -'sd65019;
    data[ 4782] =  'sd36390;
    data[ 4783] = -'sd72952;
    data[ 4784] = -'sd19141;
    data[ 4785] =  'sd29854;
    data[ 4786] =  'sd45137;
    data[ 4787] = -'sd11723;
    data[ 4788] =  'sd81780;
    data[ 4789] =  'sd80937;
    data[ 4790] =  'sd75036;
    data[ 4791] =  'sd33729;
    data[ 4792] =  'sd72262;
    data[ 4793] =  'sd14311;
    data[ 4794] = -'sd63664;
    data[ 4795] =  'sd45875;
    data[ 4796] = -'sd6557;
    data[ 4797] = -'sd45899;
    data[ 4798] =  'sd6389;
    data[ 4799] =  'sd44723;
    data[ 4800] = -'sd14621;
    data[ 4801] =  'sd61494;
    data[ 4802] = -'sd61065;
    data[ 4803] =  'sd64068;
    data[ 4804] = -'sd43047;
    data[ 4805] =  'sd26353;
    data[ 4806] =  'sd20630;
    data[ 4807] = -'sd19431;
    data[ 4808] =  'sd27824;
    data[ 4809] =  'sd30927;
    data[ 4810] =  'sd52648;
    data[ 4811] =  'sd40854;
    data[ 4812] = -'sd41704;
    data[ 4813] =  'sd35754;
    data[ 4814] = -'sd77404;
    data[ 4815] = -'sd50305;
    data[ 4816] = -'sd24453;
    data[ 4817] = -'sd7330;
    data[ 4818] = -'sd51310;
    data[ 4819] = -'sd31488;
    data[ 4820] = -'sd56575;
    data[ 4821] = -'sd68343;
    data[ 4822] =  'sd13122;
    data[ 4823] = -'sd71987;
    data[ 4824] = -'sd12386;
    data[ 4825] =  'sd77139;
    data[ 4826] =  'sd48450;
    data[ 4827] =  'sd11468;
    data[ 4828] =  'sd80276;
    data[ 4829] =  'sd70409;
    data[ 4830] =  'sd1340;
    data[ 4831] =  'sd9380;
    data[ 4832] =  'sd65660;
    data[ 4833] = -'sd31903;
    data[ 4834] = -'sd59480;
    data[ 4835] =  'sd75163;
    data[ 4836] =  'sd34618;
    data[ 4837] =  'sd78485;
    data[ 4838] =  'sd57872;
    data[ 4839] =  'sd77422;
    data[ 4840] =  'sd50431;
    data[ 4841] =  'sd25335;
    data[ 4842] =  'sd13504;
    data[ 4843] = -'sd69313;
    data[ 4844] =  'sd6332;
    data[ 4845] =  'sd44324;
    data[ 4846] = -'sd17414;
    data[ 4847] =  'sd41943;
    data[ 4848] = -'sd34081;
    data[ 4849] = -'sd74726;
    data[ 4850] = -'sd31559;
    data[ 4851] = -'sd57072;
    data[ 4852] = -'sd71822;
    data[ 4853] = -'sd11231;
    data[ 4854] = -'sd78617;
    data[ 4855] = -'sd58796;
    data[ 4856] =  'sd79951;
    data[ 4857] =  'sd68134;
    data[ 4858] = -'sd14585;
    data[ 4859] =  'sd61746;
    data[ 4860] = -'sd59301;
    data[ 4861] =  'sd76416;
    data[ 4862] =  'sd43389;
    data[ 4863] = -'sd23959;
    data[ 4864] = -'sd3872;
    data[ 4865] = -'sd27104;
    data[ 4866] = -'sd25887;
    data[ 4867] = -'sd17368;
    data[ 4868] =  'sd42265;
    data[ 4869] = -'sd31827;
    data[ 4870] = -'sd58948;
    data[ 4871] =  'sd78887;
    data[ 4872] =  'sd60686;
    data[ 4873] = -'sd66721;
    data[ 4874] =  'sd24476;
    data[ 4875] =  'sd7491;
    data[ 4876] =  'sd52437;
    data[ 4877] =  'sd39377;
    data[ 4878] = -'sd52043;
    data[ 4879] = -'sd36619;
    data[ 4880] =  'sd71349;
    data[ 4881] =  'sd7920;
    data[ 4882] =  'sd55440;
    data[ 4883] =  'sd60398;
    data[ 4884] = -'sd68737;
    data[ 4885] =  'sd10364;
    data[ 4886] =  'sd72548;
    data[ 4887] =  'sd16313;
    data[ 4888] = -'sd49650;
    data[ 4889] = -'sd19868;
    data[ 4890] =  'sd24765;
    data[ 4891] =  'sd9514;
    data[ 4892] =  'sd66598;
    data[ 4893] = -'sd25337;
    data[ 4894] = -'sd13518;
    data[ 4895] =  'sd69215;
    data[ 4896] = -'sd7018;
    data[ 4897] = -'sd49126;
    data[ 4898] = -'sd16200;
    data[ 4899] =  'sd50441;
    data[ 4900] =  'sd25405;
    data[ 4901] =  'sd13994;
    data[ 4902] = -'sd65883;
    data[ 4903] =  'sd30342;
    data[ 4904] =  'sd48553;
    data[ 4905] =  'sd12189;
    data[ 4906] = -'sd78518;
    data[ 4907] = -'sd58103;
    data[ 4908] = -'sd79039;
    data[ 4909] = -'sd61750;
    data[ 4910] =  'sd59273;
    data[ 4911] = -'sd76612;
    data[ 4912] = -'sd44761;
    data[ 4913] =  'sd14355;
    data[ 4914] = -'sd63356;
    data[ 4915] =  'sd48031;
    data[ 4916] =  'sd8535;
    data[ 4917] =  'sd59745;
    data[ 4918] = -'sd73308;
    data[ 4919] = -'sd21633;
    data[ 4920] =  'sd12410;
    data[ 4921] = -'sd76971;
    data[ 4922] = -'sd47274;
    data[ 4923] = -'sd3236;
    data[ 4924] = -'sd22652;
    data[ 4925] =  'sd5277;
    data[ 4926] =  'sd36939;
    data[ 4927] = -'sd69109;
    data[ 4928] =  'sd7760;
    data[ 4929] =  'sd54320;
    data[ 4930] =  'sd52558;
    data[ 4931] =  'sd40224;
    data[ 4932] = -'sd46114;
    data[ 4933] =  'sd4884;
    data[ 4934] =  'sd34188;
    data[ 4935] =  'sd75475;
    data[ 4936] =  'sd36802;
    data[ 4937] = -'sd70068;
    data[ 4938] =  'sd1047;
    data[ 4939] =  'sd7329;
    data[ 4940] =  'sd51303;
    data[ 4941] =  'sd31439;
    data[ 4942] =  'sd56232;
    data[ 4943] =  'sd65942;
    data[ 4944] = -'sd29929;
    data[ 4945] = -'sd45662;
    data[ 4946] =  'sd8048;
    data[ 4947] =  'sd56336;
    data[ 4948] =  'sd66670;
    data[ 4949] = -'sd24833;
    data[ 4950] = -'sd9990;
    data[ 4951] = -'sd69930;
    data[ 4952] =  'sd2013;
    data[ 4953] =  'sd14091;
    data[ 4954] = -'sd65204;
    data[ 4955] =  'sd35095;
    data[ 4956] =  'sd81824;
    data[ 4957] =  'sd81245;
    data[ 4958] =  'sd77192;
    data[ 4959] =  'sd48821;
    data[ 4960] =  'sd14065;
    data[ 4961] = -'sd65386;
    data[ 4962] =  'sd33821;
    data[ 4963] =  'sd72906;
    data[ 4964] =  'sd18819;
    data[ 4965] = -'sd32108;
    data[ 4966] = -'sd60915;
    data[ 4967] =  'sd65118;
    data[ 4968] = -'sd35697;
    data[ 4969] =  'sd77803;
    data[ 4970] =  'sd53098;
    data[ 4971] =  'sd44004;
    data[ 4972] = -'sd19654;
    data[ 4973] =  'sd26263;
    data[ 4974] =  'sd20000;
    data[ 4975] = -'sd23841;
    data[ 4976] = -'sd3046;
    data[ 4977] = -'sd21322;
    data[ 4978] =  'sd14587;
    data[ 4979] = -'sd61732;
    data[ 4980] =  'sd59399;
    data[ 4981] = -'sd75730;
    data[ 4982] = -'sd38587;
    data[ 4983] =  'sd57573;
    data[ 4984] =  'sd75329;
    data[ 4985] =  'sd35780;
    data[ 4986] = -'sd77222;
    data[ 4987] = -'sd49031;
    data[ 4988] = -'sd15535;
    data[ 4989] =  'sd55096;
    data[ 4990] =  'sd57990;
    data[ 4991] =  'sd78248;
    data[ 4992] =  'sd56213;
    data[ 4993] =  'sd65809;
    data[ 4994] = -'sd30860;
    data[ 4995] = -'sd52179;
    data[ 4996] = -'sd37571;
    data[ 4997] =  'sd64685;
    data[ 4998] = -'sd38728;
    data[ 4999] =  'sd56586;
    data[ 5000] =  'sd68420;
    data[ 5001] = -'sd12583;
    data[ 5002] =  'sd75760;
    data[ 5003] =  'sd38797;
    data[ 5004] = -'sd56103;
    data[ 5005] = -'sd65039;
    data[ 5006] =  'sd36250;
    data[ 5007] = -'sd73932;
    data[ 5008] = -'sd26001;
    data[ 5009] = -'sd18166;
    data[ 5010] =  'sd36679;
    data[ 5011] = -'sd70929;
    data[ 5012] = -'sd4980;
    data[ 5013] = -'sd34860;
    data[ 5014] = -'sd80179;
    data[ 5015] = -'sd69730;
    data[ 5016] =  'sd3413;
    data[ 5017] =  'sd23891;
    data[ 5018] =  'sd3396;
    data[ 5019] =  'sd23772;
    data[ 5020] =  'sd2563;
    data[ 5021] =  'sd17941;
    data[ 5022] = -'sd38254;
    data[ 5023] =  'sd59904;
    data[ 5024] = -'sd72195;
    data[ 5025] = -'sd13842;
    data[ 5026] =  'sd66947;
    data[ 5027] = -'sd22894;
    data[ 5028] =  'sd3583;
    data[ 5029] =  'sd25081;
    data[ 5030] =  'sd11726;
    data[ 5031] = -'sd81759;
    data[ 5032] = -'sd80790;
    data[ 5033] = -'sd74007;
    data[ 5034] = -'sd26526;
    data[ 5035] = -'sd21841;
    data[ 5036] =  'sd10954;
    data[ 5037] =  'sd76678;
    data[ 5038] =  'sd45223;
    data[ 5039] = -'sd11121;
    data[ 5040] = -'sd77847;
    data[ 5041] = -'sd53406;
    data[ 5042] = -'sd46160;
    data[ 5043] =  'sd4562;
    data[ 5044] =  'sd31934;
    data[ 5045] =  'sd59697;
    data[ 5046] = -'sd73644;
    data[ 5047] = -'sd23985;
    data[ 5048] = -'sd4054;
    data[ 5049] = -'sd28378;
    data[ 5050] = -'sd34805;
    data[ 5051] = -'sd79794;
    data[ 5052] = -'sd67035;
    data[ 5053] =  'sd22278;
    data[ 5054] = -'sd7895;
    data[ 5055] = -'sd55265;
    data[ 5056] = -'sd59173;
    data[ 5057] =  'sd77312;
    data[ 5058] =  'sd49661;
    data[ 5059] =  'sd19945;
    data[ 5060] = -'sd24226;
    data[ 5061] = -'sd5741;
    data[ 5062] = -'sd40187;
    data[ 5063] =  'sd46373;
    data[ 5064] = -'sd3071;
    data[ 5065] = -'sd21497;
    data[ 5066] =  'sd13362;
    data[ 5067] = -'sd70307;
    data[ 5068] = -'sd626;
    data[ 5069] = -'sd4382;
    data[ 5070] = -'sd30674;
    data[ 5071] = -'sd50877;
    data[ 5072] = -'sd28457;
    data[ 5073] = -'sd35358;
    data[ 5074] =  'sd80176;
    data[ 5075] =  'sd69709;
    data[ 5076] = -'sd3560;
    data[ 5077] = -'sd24920;
    data[ 5078] = -'sd10599;
    data[ 5079] = -'sd74193;
    data[ 5080] = -'sd27828;
    data[ 5081] = -'sd30955;
    data[ 5082] = -'sd52844;
    data[ 5083] = -'sd42226;
    data[ 5084] =  'sd32100;
    data[ 5085] =  'sd60859;
    data[ 5086] = -'sd65510;
    data[ 5087] =  'sd32953;
    data[ 5088] =  'sd66830;
    data[ 5089] = -'sd23713;
    data[ 5090] = -'sd2150;
    data[ 5091] = -'sd15050;
    data[ 5092] =  'sd58491;
    data[ 5093] =  'sd81755;
    data[ 5094] =  'sd80762;
    data[ 5095] =  'sd73811;
    data[ 5096] =  'sd25154;
    data[ 5097] =  'sd12237;
    data[ 5098] = -'sd78182;
    data[ 5099] = -'sd55751;
    data[ 5100] = -'sd62575;
    data[ 5101] =  'sd53498;
    data[ 5102] =  'sd46804;
    data[ 5103] = -'sd54;
    data[ 5104] = -'sd378;
    data[ 5105] = -'sd2646;
    data[ 5106] = -'sd18522;
    data[ 5107] =  'sd34187;
    data[ 5108] =  'sd75468;
    data[ 5109] =  'sd36753;
    data[ 5110] = -'sd70411;
    data[ 5111] = -'sd1354;
    data[ 5112] = -'sd9478;
    data[ 5113] = -'sd66346;
    data[ 5114] =  'sd27101;
    data[ 5115] =  'sd25866;
    data[ 5116] =  'sd17221;
    data[ 5117] = -'sd43294;
    data[ 5118] =  'sd24624;
    data[ 5119] =  'sd8527;
    data[ 5120] =  'sd59689;
    data[ 5121] = -'sd73700;
    data[ 5122] = -'sd24377;
    data[ 5123] = -'sd6798;
    data[ 5124] = -'sd47586;
    data[ 5125] = -'sd5420;
    data[ 5126] = -'sd37940;
    data[ 5127] =  'sd62102;
    data[ 5128] = -'sd56809;
    data[ 5129] = -'sd69981;
    data[ 5130] =  'sd1656;
    data[ 5131] =  'sd11592;
    data[ 5132] =  'sd81144;
    data[ 5133] =  'sd76485;
    data[ 5134] =  'sd43872;
    data[ 5135] = -'sd20578;
    data[ 5136] =  'sd19795;
    data[ 5137] = -'sd25276;
    data[ 5138] = -'sd13091;
    data[ 5139] =  'sd72204;
    data[ 5140] =  'sd13905;
    data[ 5141] = -'sd66506;
    data[ 5142] =  'sd25981;
    data[ 5143] =  'sd18026;
    data[ 5144] = -'sd37659;
    data[ 5145] =  'sd64069;
    data[ 5146] = -'sd43040;
    data[ 5147] =  'sd26402;
    data[ 5148] =  'sd20973;
    data[ 5149] = -'sd17030;
    data[ 5150] =  'sd44631;
    data[ 5151] = -'sd15265;
    data[ 5152] =  'sd56986;
    data[ 5153] =  'sd71220;
    data[ 5154] =  'sd7017;
    data[ 5155] =  'sd49119;
    data[ 5156] =  'sd16151;
    data[ 5157] = -'sd50784;
    data[ 5158] = -'sd27806;
    data[ 5159] = -'sd30801;
    data[ 5160] = -'sd51766;
    data[ 5161] = -'sd34680;
    data[ 5162] = -'sd78919;
    data[ 5163] = -'sd60910;
    data[ 5164] =  'sd65153;
    data[ 5165] = -'sd35452;
    data[ 5166] =  'sd79518;
    data[ 5167] =  'sd65103;
    data[ 5168] = -'sd35802;
    data[ 5169] =  'sd77068;
    data[ 5170] =  'sd47953;
    data[ 5171] =  'sd7989;
    data[ 5172] =  'sd55923;
    data[ 5173] =  'sd63779;
    data[ 5174] = -'sd45070;
    data[ 5175] =  'sd12192;
    data[ 5176] = -'sd78497;
    data[ 5177] = -'sd57956;
    data[ 5178] = -'sd78010;
    data[ 5179] = -'sd54547;
    data[ 5180] = -'sd54147;
    data[ 5181] = -'sd51347;
    data[ 5182] = -'sd31747;
    data[ 5183] = -'sd58388;
    data[ 5184] = -'sd81034;
    data[ 5185] = -'sd75715;
    data[ 5186] = -'sd38482;
    data[ 5187] =  'sd58308;
    data[ 5188] =  'sd80474;
    data[ 5189] =  'sd71795;
    data[ 5190] =  'sd11042;
    data[ 5191] =  'sd77294;
    data[ 5192] =  'sd49535;
    data[ 5193] =  'sd19063;
    data[ 5194] = -'sd30400;
    data[ 5195] = -'sd48959;
    data[ 5196] = -'sd15031;
    data[ 5197] =  'sd58624;
    data[ 5198] = -'sd81155;
    data[ 5199] = -'sd76562;
    data[ 5200] = -'sd44411;
    data[ 5201] =  'sd16805;
    data[ 5202] = -'sd46206;
    data[ 5203] =  'sd4240;
    data[ 5204] =  'sd29680;
    data[ 5205] =  'sd43919;
    data[ 5206] = -'sd20249;
    data[ 5207] =  'sd22098;
    data[ 5208] = -'sd9155;
    data[ 5209] = -'sd64085;
    data[ 5210] =  'sd42928;
    data[ 5211] = -'sd27186;
    data[ 5212] = -'sd26461;
    data[ 5213] = -'sd21386;
    data[ 5214] =  'sd14139;
    data[ 5215] = -'sd64868;
    data[ 5216] =  'sd37447;
    data[ 5217] = -'sd65553;
    data[ 5218] =  'sd32652;
    data[ 5219] =  'sd64723;
    data[ 5220] = -'sd38462;
    data[ 5221] =  'sd58448;
    data[ 5222] =  'sd81454;
    data[ 5223] =  'sd78655;
    data[ 5224] =  'sd59062;
    data[ 5225] = -'sd78089;
    data[ 5226] = -'sd55100;
    data[ 5227] = -'sd58018;
    data[ 5228] = -'sd78444;
    data[ 5229] = -'sd57585;
    data[ 5230] = -'sd75413;
    data[ 5231] = -'sd36368;
    data[ 5232] =  'sd73106;
    data[ 5233] =  'sd20219;
    data[ 5234] = -'sd22308;
    data[ 5235] =  'sd7685;
    data[ 5236] =  'sd53795;
    data[ 5237] =  'sd48883;
    data[ 5238] =  'sd14499;
    data[ 5239] = -'sd62348;
    data[ 5240] =  'sd55087;
    data[ 5241] =  'sd57927;
    data[ 5242] =  'sd77807;
    data[ 5243] =  'sd53126;
    data[ 5244] =  'sd44200;
    data[ 5245] = -'sd18282;
    data[ 5246] =  'sd35867;
    data[ 5247] = -'sd76613;
    data[ 5248] = -'sd44768;
    data[ 5249] =  'sd14306;
    data[ 5250] = -'sd63699;
    data[ 5251] =  'sd45630;
    data[ 5252] = -'sd8272;
    data[ 5253] = -'sd57904;
    data[ 5254] = -'sd77646;
    data[ 5255] = -'sd51999;
    data[ 5256] = -'sd36311;
    data[ 5257] =  'sd73505;
    data[ 5258] =  'sd23012;
    data[ 5259] = -'sd2757;
    data[ 5260] = -'sd19299;
    data[ 5261] =  'sd28748;
    data[ 5262] =  'sd37395;
    data[ 5263] = -'sd65917;
    data[ 5264] =  'sd30104;
    data[ 5265] =  'sd46887;
    data[ 5266] =  'sd527;
    data[ 5267] =  'sd3689;
    data[ 5268] =  'sd25823;
    data[ 5269] =  'sd16920;
    data[ 5270] = -'sd45401;
    data[ 5271] =  'sd9875;
    data[ 5272] =  'sd69125;
    data[ 5273] = -'sd7648;
    data[ 5274] = -'sd53536;
    data[ 5275] = -'sd47070;
    data[ 5276] = -'sd1808;
    data[ 5277] = -'sd12656;
    data[ 5278] =  'sd75249;
    data[ 5279] =  'sd35220;
    data[ 5280] = -'sd81142;
    data[ 5281] = -'sd76471;
    data[ 5282] = -'sd43774;
    data[ 5283] =  'sd21264;
    data[ 5284] = -'sd14993;
    data[ 5285] =  'sd58890;
    data[ 5286] = -'sd79293;
    data[ 5287] = -'sd63528;
    data[ 5288] =  'sd46827;
    data[ 5289] =  'sd107;
    data[ 5290] =  'sd749;
    data[ 5291] =  'sd5243;
    data[ 5292] =  'sd36701;
    data[ 5293] = -'sd70775;
    data[ 5294] = -'sd3902;
    data[ 5295] = -'sd27314;
    data[ 5296] = -'sd27357;
    data[ 5297] = -'sd27658;
    data[ 5298] = -'sd29765;
    data[ 5299] = -'sd44514;
    data[ 5300] =  'sd16084;
    data[ 5301] = -'sd51253;
    data[ 5302] = -'sd31089;
    data[ 5303] = -'sd53782;
    data[ 5304] = -'sd48792;
    data[ 5305] = -'sd13862;
    data[ 5306] =  'sd66807;
    data[ 5307] = -'sd23874;
    data[ 5308] = -'sd3277;
    data[ 5309] = -'sd22939;
    data[ 5310] =  'sd3268;
    data[ 5311] =  'sd22876;
    data[ 5312] = -'sd3709;
    data[ 5313] = -'sd25963;
    data[ 5314] = -'sd17900;
    data[ 5315] =  'sd38541;
    data[ 5316] = -'sd57895;
    data[ 5317] = -'sd77583;
    data[ 5318] = -'sd51558;
    data[ 5319] = -'sd33224;
    data[ 5320] = -'sd68727;
    data[ 5321] =  'sd10434;
    data[ 5322] =  'sd73038;
    data[ 5323] =  'sd19743;
    data[ 5324] = -'sd25640;
    data[ 5325] = -'sd15639;
    data[ 5326] =  'sd54368;
    data[ 5327] =  'sd52894;
    data[ 5328] =  'sd42576;
    data[ 5329] = -'sd29650;
    data[ 5330] = -'sd43709;
    data[ 5331] =  'sd21719;
    data[ 5332] = -'sd11808;
    data[ 5333] =  'sd81185;
    data[ 5334] =  'sd76772;
    data[ 5335] =  'sd45881;
    data[ 5336] = -'sd6515;
    data[ 5337] = -'sd45605;
    data[ 5338] =  'sd8447;
    data[ 5339] =  'sd59129;
    data[ 5340] = -'sd77620;
    data[ 5341] = -'sd51817;
    data[ 5342] = -'sd35037;
    data[ 5343] = -'sd81418;
    data[ 5344] = -'sd78403;
    data[ 5345] = -'sd57298;
    data[ 5346] = -'sd73404;
    data[ 5347] = -'sd22305;
    data[ 5348] =  'sd7706;
    data[ 5349] =  'sd53942;
    data[ 5350] =  'sd49912;
    data[ 5351] =  'sd21702;
    data[ 5352] = -'sd11927;
    data[ 5353] =  'sd80352;
    data[ 5354] =  'sd70941;
    data[ 5355] =  'sd5064;
    data[ 5356] =  'sd35448;
    data[ 5357] = -'sd79546;
    data[ 5358] = -'sd65299;
    data[ 5359] =  'sd34430;
    data[ 5360] =  'sd77169;
    data[ 5361] =  'sd48660;
    data[ 5362] =  'sd12938;
    data[ 5363] = -'sd73275;
    data[ 5364] = -'sd21402;
    data[ 5365] =  'sd14027;
    data[ 5366] = -'sd65652;
    data[ 5367] =  'sd31959;
    data[ 5368] =  'sd59872;
    data[ 5369] = -'sd72419;
    data[ 5370] = -'sd15410;
    data[ 5371] =  'sd55971;
    data[ 5372] =  'sd64115;
    data[ 5373] = -'sd42718;
    data[ 5374] =  'sd28656;
    data[ 5375] =  'sd36751;
    data[ 5376] = -'sd70425;
    data[ 5377] = -'sd1452;
    data[ 5378] = -'sd10164;
    data[ 5379] = -'sd71148;
    data[ 5380] = -'sd6513;
    data[ 5381] = -'sd45591;
    data[ 5382] =  'sd8545;
    data[ 5383] =  'sd59815;
    data[ 5384] = -'sd72818;
    data[ 5385] = -'sd18203;
    data[ 5386] =  'sd36420;
    data[ 5387] = -'sd72742;
    data[ 5388] = -'sd17671;
    data[ 5389] =  'sd40144;
    data[ 5390] = -'sd46674;
    data[ 5391] =  'sd964;
    data[ 5392] =  'sd6748;
    data[ 5393] =  'sd47236;
    data[ 5394] =  'sd2970;
    data[ 5395] =  'sd20790;
    data[ 5396] = -'sd18311;
    data[ 5397] =  'sd35664;
    data[ 5398] = -'sd78034;
    data[ 5399] = -'sd54715;
    data[ 5400] = -'sd55323;
    data[ 5401] = -'sd59579;
    data[ 5402] =  'sd74470;
    data[ 5403] =  'sd29767;
    data[ 5404] =  'sd44528;
    data[ 5405] = -'sd15986;
    data[ 5406] =  'sd51939;
    data[ 5407] =  'sd35891;
    data[ 5408] = -'sd76445;
    data[ 5409] = -'sd43592;
    data[ 5410] =  'sd22538;
    data[ 5411] = -'sd6075;
    data[ 5412] = -'sd42525;
    data[ 5413] =  'sd30007;
    data[ 5414] =  'sd46208;
    data[ 5415] = -'sd4226;
    data[ 5416] = -'sd29582;
    data[ 5417] = -'sd43233;
    data[ 5418] =  'sd25051;
    data[ 5419] =  'sd11516;
    data[ 5420] =  'sd80612;
    data[ 5421] =  'sd72761;
    data[ 5422] =  'sd17804;
    data[ 5423] = -'sd39213;
    data[ 5424] =  'sd53191;
    data[ 5425] =  'sd44655;
    data[ 5426] = -'sd15097;
    data[ 5427] =  'sd58162;
    data[ 5428] =  'sd79452;
    data[ 5429] =  'sd64641;
    data[ 5430] = -'sd39036;
    data[ 5431] =  'sd54430;
    data[ 5432] =  'sd53328;
    data[ 5433] =  'sd45614;
    data[ 5434] = -'sd8384;
    data[ 5435] = -'sd58688;
    data[ 5436] =  'sd80707;
    data[ 5437] =  'sd73426;
    data[ 5438] =  'sd22459;
    data[ 5439] = -'sd6628;
    data[ 5440] = -'sd46396;
    data[ 5441] =  'sd2910;
    data[ 5442] =  'sd20370;
    data[ 5443] = -'sd21251;
    data[ 5444] =  'sd15084;
    data[ 5445] = -'sd58253;
    data[ 5446] = -'sd80089;
    data[ 5447] = -'sd69100;
    data[ 5448] =  'sd7823;
    data[ 5449] =  'sd54761;
    data[ 5450] =  'sd55645;
    data[ 5451] =  'sd61833;
    data[ 5452] = -'sd58692;
    data[ 5453] =  'sd80679;
    data[ 5454] =  'sd73230;
    data[ 5455] =  'sd21087;
    data[ 5456] = -'sd16232;
    data[ 5457] =  'sd50217;
    data[ 5458] =  'sd23837;
    data[ 5459] =  'sd3018;
    data[ 5460] =  'sd21126;
    data[ 5461] = -'sd15959;
    data[ 5462] =  'sd52128;
    data[ 5463] =  'sd37214;
    data[ 5464] = -'sd67184;
    data[ 5465] =  'sd21235;
    data[ 5466] = -'sd15196;
    data[ 5467] =  'sd57469;
    data[ 5468] =  'sd74601;
    data[ 5469] =  'sd30684;
    data[ 5470] =  'sd50947;
    data[ 5471] =  'sd28947;
    data[ 5472] =  'sd38788;
    data[ 5473] = -'sd56166;
    data[ 5474] = -'sd65480;
    data[ 5475] =  'sd33163;
    data[ 5476] =  'sd68300;
    data[ 5477] = -'sd13423;
    data[ 5478] =  'sd69880;
    data[ 5479] = -'sd2363;
    data[ 5480] = -'sd16541;
    data[ 5481] =  'sd48054;
    data[ 5482] =  'sd8696;
    data[ 5483] =  'sd60872;
    data[ 5484] = -'sd65419;
    data[ 5485] =  'sd33590;
    data[ 5486] =  'sd71289;
    data[ 5487] =  'sd7500;
    data[ 5488] =  'sd52500;
    data[ 5489] =  'sd39818;
    data[ 5490] = -'sd48956;
    data[ 5491] = -'sd15010;
    data[ 5492] =  'sd58771;
    data[ 5493] = -'sd80126;
    data[ 5494] = -'sd69359;
    data[ 5495] =  'sd6010;
    data[ 5496] =  'sd42070;
    data[ 5497] = -'sd33192;
    data[ 5498] = -'sd68503;
    data[ 5499] =  'sd12002;
    data[ 5500] = -'sd79827;
    data[ 5501] = -'sd67266;
    data[ 5502] =  'sd20661;
    data[ 5503] = -'sd19214;
    data[ 5504] =  'sd29343;
    data[ 5505] =  'sd41560;
    data[ 5506] = -'sd36762;
    data[ 5507] =  'sd70348;
    data[ 5508] =  'sd913;
    data[ 5509] =  'sd6391;
    data[ 5510] =  'sd44737;
    data[ 5511] = -'sd14523;
    data[ 5512] =  'sd62180;
    data[ 5513] = -'sd56263;
    data[ 5514] = -'sd66159;
    data[ 5515] =  'sd28410;
    data[ 5516] =  'sd35029;
    data[ 5517] =  'sd81362;
    data[ 5518] =  'sd78011;
    data[ 5519] =  'sd54554;
    data[ 5520] =  'sd54196;
    data[ 5521] =  'sd51690;
    data[ 5522] =  'sd34148;
    data[ 5523] =  'sd75195;
    data[ 5524] =  'sd34842;
    data[ 5525] =  'sd80053;
    data[ 5526] =  'sd68848;
    data[ 5527] = -'sd9587;
    data[ 5528] = -'sd67109;
    data[ 5529] =  'sd21760;
    data[ 5530] = -'sd11521;
    data[ 5531] = -'sd80647;
    data[ 5532] = -'sd73006;
    data[ 5533] = -'sd19519;
    data[ 5534] =  'sd27208;
    data[ 5535] =  'sd26615;
    data[ 5536] =  'sd22464;
    data[ 5537] = -'sd6593;
    data[ 5538] = -'sd46151;
    data[ 5539] =  'sd4625;
    data[ 5540] =  'sd32375;
    data[ 5541] =  'sd62784;
    data[ 5542] = -'sd52035;
    data[ 5543] = -'sd36563;
    data[ 5544] =  'sd71741;
    data[ 5545] =  'sd10664;
    data[ 5546] =  'sd74648;
    data[ 5547] =  'sd31013;
    data[ 5548] =  'sd53250;
    data[ 5549] =  'sd45068;
    data[ 5550] = -'sd12206;
    data[ 5551] =  'sd78399;
    data[ 5552] =  'sd57270;
    data[ 5553] =  'sd73208;
    data[ 5554] =  'sd20933;
    data[ 5555] = -'sd17310;
    data[ 5556] =  'sd42671;
    data[ 5557] = -'sd28985;
    data[ 5558] = -'sd39054;
    data[ 5559] =  'sd54304;
    data[ 5560] =  'sd52446;
    data[ 5561] =  'sd39440;
    data[ 5562] = -'sd51602;
    data[ 5563] = -'sd33532;
    data[ 5564] = -'sd70883;
    data[ 5565] = -'sd4658;
    data[ 5566] = -'sd32606;
    data[ 5567] = -'sd64401;
    data[ 5568] =  'sd40716;
    data[ 5569] = -'sd42670;
    data[ 5570] =  'sd28992;
    data[ 5571] =  'sd39103;
    data[ 5572] = -'sd53961;
    data[ 5573] = -'sd50045;
    data[ 5574] = -'sd22633;
    data[ 5575] =  'sd5410;
    data[ 5576] =  'sd37870;
    data[ 5577] = -'sd62592;
    data[ 5578] =  'sd53379;
    data[ 5579] =  'sd45971;
    data[ 5580] = -'sd5885;
    data[ 5581] = -'sd41195;
    data[ 5582] =  'sd39317;
    data[ 5583] = -'sd52463;
    data[ 5584] = -'sd39559;
    data[ 5585] =  'sd50769;
    data[ 5586] =  'sd27701;
    data[ 5587] =  'sd30066;
    data[ 5588] =  'sd46621;
    data[ 5589] = -'sd1335;
    data[ 5590] = -'sd9345;
    data[ 5591] = -'sd65415;
    data[ 5592] =  'sd33618;
    data[ 5593] =  'sd71485;
    data[ 5594] =  'sd8872;
    data[ 5595] =  'sd62104;
    data[ 5596] = -'sd56795;
    data[ 5597] = -'sd69883;
    data[ 5598] =  'sd2342;
    data[ 5599] =  'sd16394;
    data[ 5600] = -'sd49083;
    data[ 5601] = -'sd15899;
    data[ 5602] =  'sd52548;
    data[ 5603] =  'sd40154;
    data[ 5604] = -'sd46604;
    data[ 5605] =  'sd1454;
    data[ 5606] =  'sd10178;
    data[ 5607] =  'sd71246;
    data[ 5608] =  'sd7199;
    data[ 5609] =  'sd50393;
    data[ 5610] =  'sd25069;
    data[ 5611] =  'sd11642;
    data[ 5612] =  'sd81494;
    data[ 5613] =  'sd78935;
    data[ 5614] =  'sd61022;
    data[ 5615] = -'sd64369;
    data[ 5616] =  'sd40940;
    data[ 5617] = -'sd41102;
    data[ 5618] =  'sd39968;
    data[ 5619] = -'sd47906;
    data[ 5620] = -'sd7660;
    data[ 5621] = -'sd53620;
    data[ 5622] = -'sd47658;
    data[ 5623] = -'sd5924;
    data[ 5624] = -'sd41468;
    data[ 5625] =  'sd37406;
    data[ 5626] = -'sd65840;
    data[ 5627] =  'sd30643;
    data[ 5628] =  'sd50660;
    data[ 5629] =  'sd26938;
    data[ 5630] =  'sd24725;
    data[ 5631] =  'sd9234;
    data[ 5632] =  'sd64638;
    data[ 5633] = -'sd39057;
    data[ 5634] =  'sd54283;
    data[ 5635] =  'sd52299;
    data[ 5636] =  'sd38411;
    data[ 5637] = -'sd58805;
    data[ 5638] =  'sd79888;
    data[ 5639] =  'sd67693;
    data[ 5640] = -'sd17672;
    data[ 5641] =  'sd40137;
    data[ 5642] = -'sd46723;
    data[ 5643] =  'sd621;
    data[ 5644] =  'sd4347;
    data[ 5645] =  'sd30429;
    data[ 5646] =  'sd49162;
    data[ 5647] =  'sd16452;
    data[ 5648] = -'sd48677;
    data[ 5649] = -'sd13057;
    data[ 5650] =  'sd72442;
    data[ 5651] =  'sd15571;
    data[ 5652] = -'sd54844;
    data[ 5653] = -'sd56226;
    data[ 5654] = -'sd65900;
    data[ 5655] =  'sd30223;
    data[ 5656] =  'sd47720;
    data[ 5657] =  'sd6358;
    data[ 5658] =  'sd44506;
    data[ 5659] = -'sd16140;
    data[ 5660] =  'sd50861;
    data[ 5661] =  'sd28345;
    data[ 5662] =  'sd34574;
    data[ 5663] =  'sd78177;
    data[ 5664] =  'sd55716;
    data[ 5665] =  'sd62330;
    data[ 5666] = -'sd55213;
    data[ 5667] = -'sd58809;
    data[ 5668] =  'sd79860;
    data[ 5669] =  'sd67497;
    data[ 5670] = -'sd19044;
    data[ 5671] =  'sd30533;
    data[ 5672] =  'sd49890;
    data[ 5673] =  'sd21548;
    data[ 5674] = -'sd13005;
    data[ 5675] =  'sd72806;
    data[ 5676] =  'sd18119;
    data[ 5677] = -'sd37008;
    data[ 5678] =  'sd68626;
    data[ 5679] = -'sd11141;
    data[ 5680] = -'sd77987;
    data[ 5681] = -'sd54386;
    data[ 5682] = -'sd53020;
    data[ 5683] = -'sd43458;
    data[ 5684] =  'sd23476;
    data[ 5685] =  'sd491;
    data[ 5686] =  'sd3437;
    data[ 5687] =  'sd24059;
    data[ 5688] =  'sd4572;
    data[ 5689] =  'sd32004;
    data[ 5690] =  'sd60187;
    data[ 5691] = -'sd70214;
    data[ 5692] =  'sd25;
    data[ 5693] =  'sd175;
    data[ 5694] =  'sd1225;
    data[ 5695] =  'sd8575;
    data[ 5696] =  'sd60025;
    data[ 5697] = -'sd71348;
    data[ 5698] = -'sd7913;
    data[ 5699] = -'sd55391;
    data[ 5700] = -'sd60055;
    data[ 5701] =  'sd71138;
    data[ 5702] =  'sd6443;
    data[ 5703] =  'sd45101;
    data[ 5704] = -'sd11975;
    data[ 5705] =  'sd80016;
    data[ 5706] =  'sd68589;
    data[ 5707] = -'sd11400;
    data[ 5708] = -'sd79800;
    data[ 5709] = -'sd67077;
    data[ 5710] =  'sd21984;
    data[ 5711] = -'sd9953;
    data[ 5712] = -'sd69671;
    data[ 5713] =  'sd3826;
    data[ 5714] =  'sd26782;
    data[ 5715] =  'sd23633;
    data[ 5716] =  'sd1590;
    data[ 5717] =  'sd11130;
    data[ 5718] =  'sd77910;
    data[ 5719] =  'sd53847;
    data[ 5720] =  'sd49247;
    data[ 5721] =  'sd17047;
    data[ 5722] = -'sd44512;
    data[ 5723] =  'sd16098;
    data[ 5724] = -'sd51155;
    data[ 5725] = -'sd30403;
    data[ 5726] = -'sd48980;
    data[ 5727] = -'sd15178;
    data[ 5728] =  'sd57595;
    data[ 5729] =  'sd75483;
    data[ 5730] =  'sd36858;
    data[ 5731] = -'sd69676;
    data[ 5732] =  'sd3791;
    data[ 5733] =  'sd26537;
    data[ 5734] =  'sd21918;
    data[ 5735] = -'sd10415;
    data[ 5736] = -'sd72905;
    data[ 5737] = -'sd18812;
    data[ 5738] =  'sd32157;
    data[ 5739] =  'sd61258;
    data[ 5740] = -'sd62717;
    data[ 5741] =  'sd52504;
    data[ 5742] =  'sd39846;
    data[ 5743] = -'sd48760;
    data[ 5744] = -'sd13638;
    data[ 5745] =  'sd68375;
    data[ 5746] = -'sd12898;
    data[ 5747] =  'sd73555;
    data[ 5748] =  'sd23362;
    data[ 5749] = -'sd307;
    data[ 5750] = -'sd2149;
    data[ 5751] = -'sd15043;
    data[ 5752] =  'sd58540;
    data[ 5753] = -'sd81743;
    data[ 5754] = -'sd80678;
    data[ 5755] = -'sd73223;
    data[ 5756] = -'sd21038;
    data[ 5757] =  'sd16575;
    data[ 5758] = -'sd47816;
    data[ 5759] = -'sd7030;
    data[ 5760] = -'sd49210;
    data[ 5761] = -'sd16788;
    data[ 5762] =  'sd46325;
    data[ 5763] = -'sd3407;
    data[ 5764] = -'sd23849;
    data[ 5765] = -'sd3102;
    data[ 5766] = -'sd21714;
    data[ 5767] =  'sd11843;
    data[ 5768] = -'sd80940;
    data[ 5769] = -'sd75057;
    data[ 5770] = -'sd33876;
    data[ 5771] = -'sd73291;
    data[ 5772] = -'sd21514;
    data[ 5773] =  'sd13243;
    data[ 5774] = -'sd71140;
    data[ 5775] = -'sd6457;
    data[ 5776] = -'sd45199;
    data[ 5777] =  'sd11289;
    data[ 5778] =  'sd79023;
    data[ 5779] =  'sd61638;
    data[ 5780] = -'sd60057;
    data[ 5781] =  'sd71124;
    data[ 5782] =  'sd6345;
    data[ 5783] =  'sd44415;
    data[ 5784] = -'sd16777;
    data[ 5785] =  'sd46402;
    data[ 5786] = -'sd2868;
    data[ 5787] = -'sd20076;
    data[ 5788] =  'sd23309;
    data[ 5789] = -'sd678;
    data[ 5790] = -'sd4746;
    data[ 5791] = -'sd33222;
    data[ 5792] = -'sd68713;
    data[ 5793] =  'sd10532;
    data[ 5794] =  'sd73724;
    data[ 5795] =  'sd24545;
    data[ 5796] =  'sd7974;
    data[ 5797] =  'sd55818;
    data[ 5798] =  'sd63044;
    data[ 5799] = -'sd50215;
    data[ 5800] = -'sd23823;
    data[ 5801] = -'sd2920;
    data[ 5802] = -'sd20440;
    data[ 5803] =  'sd20761;
    data[ 5804] = -'sd18514;
    data[ 5805] =  'sd34243;
    data[ 5806] =  'sd75860;
    data[ 5807] =  'sd39497;
    data[ 5808] = -'sd51203;
    data[ 5809] = -'sd30739;
    data[ 5810] = -'sd51332;
    data[ 5811] = -'sd31642;
    data[ 5812] = -'sd57653;
    data[ 5813] = -'sd75889;
    data[ 5814] = -'sd39700;
    data[ 5815] =  'sd49782;
    data[ 5816] =  'sd20792;
    data[ 5817] = -'sd18297;
    data[ 5818] =  'sd35762;
    data[ 5819] = -'sd77348;
    data[ 5820] = -'sd49913;
    data[ 5821] = -'sd21709;
    data[ 5822] =  'sd11878;
    data[ 5823] = -'sd80695;
    data[ 5824] = -'sd73342;
    data[ 5825] = -'sd21871;
    data[ 5826] =  'sd10744;
    data[ 5827] =  'sd75208;
    data[ 5828] =  'sd34933;
    data[ 5829] =  'sd80690;
    data[ 5830] =  'sd73307;
    data[ 5831] =  'sd21626;
    data[ 5832] = -'sd12459;
    data[ 5833] =  'sd76628;
    data[ 5834] =  'sd44873;
    data[ 5835] = -'sd13571;
    data[ 5836] =  'sd68844;
    data[ 5837] = -'sd9615;
    data[ 5838] = -'sd67305;
    data[ 5839] =  'sd20388;
    data[ 5840] = -'sd21125;
    data[ 5841] =  'sd15966;
    data[ 5842] = -'sd52079;
    data[ 5843] = -'sd36871;
    data[ 5844] =  'sd69585;
    data[ 5845] = -'sd4428;
    data[ 5846] = -'sd30996;
    data[ 5847] = -'sd53131;
    data[ 5848] = -'sd44235;
    data[ 5849] =  'sd18037;
    data[ 5850] = -'sd37582;
    data[ 5851] =  'sd64608;
    data[ 5852] = -'sd39267;
    data[ 5853] =  'sd52813;
    data[ 5854] =  'sd42009;
    data[ 5855] = -'sd33619;
    data[ 5856] = -'sd71492;
    data[ 5857] = -'sd8921;
    data[ 5858] = -'sd62447;
    data[ 5859] =  'sd54394;
    data[ 5860] =  'sd53076;
    data[ 5861] =  'sd43850;
    data[ 5862] = -'sd20732;
    data[ 5863] =  'sd18717;
    data[ 5864] = -'sd32822;
    data[ 5865] = -'sd65913;
    data[ 5866] =  'sd30132;
    data[ 5867] =  'sd47083;
    data[ 5868] =  'sd1899;
    data[ 5869] =  'sd13293;
    data[ 5870] = -'sd70790;
    data[ 5871] = -'sd4007;
    data[ 5872] = -'sd28049;
    data[ 5873] = -'sd32502;
    data[ 5874] = -'sd63673;
    data[ 5875] =  'sd45812;
    data[ 5876] = -'sd6998;
    data[ 5877] = -'sd48986;
    data[ 5878] = -'sd15220;
    data[ 5879] =  'sd57301;
    data[ 5880] =  'sd73425;
    data[ 5881] =  'sd22452;
    data[ 5882] = -'sd6677;
    data[ 5883] = -'sd46739;
    data[ 5884] =  'sd509;
    data[ 5885] =  'sd3563;
    data[ 5886] =  'sd24941;
    data[ 5887] =  'sd10746;
    data[ 5888] =  'sd75222;
    data[ 5889] =  'sd35031;
    data[ 5890] =  'sd81376;
    data[ 5891] =  'sd78109;
    data[ 5892] =  'sd55240;
    data[ 5893] =  'sd58998;
    data[ 5894] = -'sd78537;
    data[ 5895] = -'sd58236;
    data[ 5896] = -'sd79970;
    data[ 5897] = -'sd68267;
    data[ 5898] =  'sd13654;
    data[ 5899] = -'sd68263;
    data[ 5900] =  'sd13682;
    data[ 5901] = -'sd68067;
    data[ 5902] =  'sd15054;
    data[ 5903] = -'sd58463;
    data[ 5904] = -'sd81559;
    data[ 5905] = -'sd79390;
    data[ 5906] = -'sd64207;
    data[ 5907] =  'sd42074;
    data[ 5908] = -'sd33164;
    data[ 5909] = -'sd68307;
    data[ 5910] =  'sd13374;
    data[ 5911] = -'sd70223;
    data[ 5912] = -'sd38;
    data[ 5913] = -'sd266;
    data[ 5914] = -'sd1862;
    data[ 5915] = -'sd13034;
    data[ 5916] =  'sd72603;
    data[ 5917] =  'sd16698;
    data[ 5918] = -'sd46955;
    data[ 5919] = -'sd1003;
    data[ 5920] = -'sd7021;
    data[ 5921] = -'sd49147;
    data[ 5922] = -'sd16347;
    data[ 5923] =  'sd49412;
    data[ 5924] =  'sd18202;
    data[ 5925] = -'sd36427;
    data[ 5926] =  'sd72693;
    data[ 5927] =  'sd17328;
    data[ 5928] = -'sd42545;
    data[ 5929] =  'sd29867;
    data[ 5930] =  'sd45228;
    data[ 5931] = -'sd11086;
    data[ 5932] = -'sd77602;
    data[ 5933] = -'sd51691;
    data[ 5934] = -'sd34155;
    data[ 5935] = -'sd75244;
    data[ 5936] = -'sd35185;
    data[ 5937] =  'sd81387;
    data[ 5938] =  'sd78186;
    data[ 5939] =  'sd55779;
    data[ 5940] =  'sd62771;
    data[ 5941] = -'sd52126;
    data[ 5942] = -'sd37200;
    data[ 5943] =  'sd67282;
    data[ 5944] = -'sd20549;
    data[ 5945] =  'sd19998;
    data[ 5946] = -'sd23855;
    data[ 5947] = -'sd3144;
    data[ 5948] = -'sd22008;
    data[ 5949] =  'sd9785;
    data[ 5950] =  'sd68495;
    data[ 5951] = -'sd12058;
    data[ 5952] =  'sd79435;
    data[ 5953] =  'sd64522;
    data[ 5954] = -'sd39869;
    data[ 5955] =  'sd48599;
    data[ 5956] =  'sd12511;
    data[ 5957] = -'sd76264;
    data[ 5958] = -'sd42325;
    data[ 5959] =  'sd31407;
    data[ 5960] =  'sd56008;
    data[ 5961] =  'sd64374;
    data[ 5962] = -'sd40905;
    data[ 5963] =  'sd41347;
    data[ 5964] = -'sd38253;
    data[ 5965] =  'sd59911;
    data[ 5966] = -'sd72146;
    data[ 5967] = -'sd13499;
    data[ 5968] =  'sd69348;
    data[ 5969] = -'sd6087;
    data[ 5970] = -'sd42609;
    data[ 5971] =  'sd29419;
    data[ 5972] =  'sd42092;
    data[ 5973] = -'sd33038;
    data[ 5974] = -'sd67425;
    data[ 5975] =  'sd19548;
    data[ 5976] = -'sd27005;
    data[ 5977] = -'sd25194;
    data[ 5978] = -'sd12517;
    data[ 5979] =  'sd76222;
    data[ 5980] =  'sd42031;
    data[ 5981] = -'sd33465;
    data[ 5982] = -'sd70414;
    data[ 5983] = -'sd1375;
    data[ 5984] = -'sd9625;
    data[ 5985] = -'sd67375;
    data[ 5986] =  'sd19898;
    data[ 5987] = -'sd24555;
    data[ 5988] = -'sd8044;
    data[ 5989] = -'sd56308;
    data[ 5990] = -'sd66474;
    data[ 5991] =  'sd26205;
    data[ 5992] =  'sd19594;
    data[ 5993] = -'sd26683;
    data[ 5994] = -'sd22940;
    data[ 5995] =  'sd3261;
    data[ 5996] =  'sd22827;
    data[ 5997] = -'sd4052;
    data[ 5998] = -'sd28364;
    data[ 5999] = -'sd34707;
    data[ 6000] = -'sd79108;
    data[ 6001] = -'sd62233;
    data[ 6002] =  'sd55892;
    data[ 6003] =  'sd63562;
    data[ 6004] = -'sd46589;
    data[ 6005] =  'sd1559;
    data[ 6006] =  'sd10913;
    data[ 6007] =  'sd76391;
    data[ 6008] =  'sd43214;
    data[ 6009] = -'sd25184;
    data[ 6010] = -'sd12447;
    data[ 6011] =  'sd76712;
    data[ 6012] =  'sd45461;
    data[ 6013] = -'sd9455;
    data[ 6014] = -'sd66185;
    data[ 6015] =  'sd28228;
    data[ 6016] =  'sd33755;
    data[ 6017] =  'sd72444;
    data[ 6018] =  'sd15585;
    data[ 6019] = -'sd54746;
    data[ 6020] = -'sd55540;
    data[ 6021] = -'sd61098;
    data[ 6022] =  'sd63837;
    data[ 6023] = -'sd44664;
    data[ 6024] =  'sd15034;
    data[ 6025] = -'sd58603;
    data[ 6026] =  'sd81302;
    data[ 6027] =  'sd77591;
    data[ 6028] =  'sd51614;
    data[ 6029] =  'sd33616;
    data[ 6030] =  'sd71471;
    data[ 6031] =  'sd8774;
    data[ 6032] =  'sd61418;
    data[ 6033] = -'sd61597;
    data[ 6034] =  'sd60344;
    data[ 6035] = -'sd69115;
    data[ 6036] =  'sd7718;
    data[ 6037] =  'sd54026;
    data[ 6038] =  'sd50500;
    data[ 6039] =  'sd25818;
    data[ 6040] =  'sd16885;
    data[ 6041] = -'sd45646;
    data[ 6042] =  'sd8160;
    data[ 6043] =  'sd57120;
    data[ 6044] =  'sd72158;
    data[ 6045] =  'sd13583;
    data[ 6046] = -'sd68760;
    data[ 6047] =  'sd10203;
    data[ 6048] =  'sd71421;
    data[ 6049] =  'sd8424;
    data[ 6050] =  'sd58968;
    data[ 6051] = -'sd78747;
    data[ 6052] = -'sd59706;
    data[ 6053] =  'sd73581;
    data[ 6054] =  'sd23544;
    data[ 6055] =  'sd967;
    data[ 6056] =  'sd6769;
    data[ 6057] =  'sd47383;
    data[ 6058] =  'sd3999;
    data[ 6059] =  'sd27993;
    data[ 6060] =  'sd32110;
    data[ 6061] =  'sd60929;
    data[ 6062] = -'sd65020;
    data[ 6063] =  'sd36383;
    data[ 6064] = -'sd73001;
    data[ 6065] = -'sd19484;
    data[ 6066] =  'sd27453;
    data[ 6067] =  'sd28330;
    data[ 6068] =  'sd34469;
    data[ 6069] =  'sd77442;
    data[ 6070] =  'sd50571;
    data[ 6071] =  'sd26315;
    data[ 6072] =  'sd20364;
    data[ 6073] = -'sd21293;
    data[ 6074] =  'sd14790;
    data[ 6075] = -'sd60311;
    data[ 6076] =  'sd69346;
    data[ 6077] = -'sd6101;
    data[ 6078] = -'sd42707;
    data[ 6079] =  'sd28733;
    data[ 6080] =  'sd37290;
    data[ 6081] = -'sd66652;
    data[ 6082] =  'sd24959;
    data[ 6083] =  'sd10872;
    data[ 6084] =  'sd76104;
    data[ 6085] =  'sd41205;
    data[ 6086] = -'sd39247;
    data[ 6087] =  'sd52953;
    data[ 6088] =  'sd42989;
    data[ 6089] = -'sd26759;
    data[ 6090] = -'sd23472;
    data[ 6091] = -'sd463;
    data[ 6092] = -'sd3241;
    data[ 6093] = -'sd22687;
    data[ 6094] =  'sd5032;
    data[ 6095] =  'sd35224;
    data[ 6096] = -'sd81114;
    data[ 6097] = -'sd76275;
    data[ 6098] = -'sd42402;
    data[ 6099] =  'sd30868;
    data[ 6100] =  'sd52235;
    data[ 6101] =  'sd37963;
    data[ 6102] = -'sd61941;
    data[ 6103] =  'sd57936;
    data[ 6104] =  'sd77870;
    data[ 6105] =  'sd53567;
    data[ 6106] =  'sd47287;
    data[ 6107] =  'sd3327;
    data[ 6108] =  'sd23289;
    data[ 6109] = -'sd818;
    data[ 6110] = -'sd5726;
    data[ 6111] = -'sd40082;
    data[ 6112] =  'sd47108;
    data[ 6113] =  'sd2074;
    data[ 6114] =  'sd14518;
    data[ 6115] = -'sd62215;
    data[ 6116] =  'sd56018;
    data[ 6117] =  'sd64444;
    data[ 6118] = -'sd40415;
    data[ 6119] =  'sd44777;
    data[ 6120] = -'sd14243;
    data[ 6121] =  'sd64140;
    data[ 6122] = -'sd42543;
    data[ 6123] =  'sd29881;
    data[ 6124] =  'sd45326;
    data[ 6125] = -'sd10400;
    data[ 6126] = -'sd72800;
    data[ 6127] = -'sd18077;
    data[ 6128] =  'sd37302;
    data[ 6129] = -'sd66568;
    data[ 6130] =  'sd25547;
    data[ 6131] =  'sd14988;
    data[ 6132] = -'sd58925;
    data[ 6133] =  'sd79048;
    data[ 6134] =  'sd61813;
    data[ 6135] = -'sd58832;
    data[ 6136] =  'sd79699;
    data[ 6137] =  'sd66370;
    data[ 6138] = -'sd26933;
    data[ 6139] = -'sd24690;
    data[ 6140] = -'sd8989;
    data[ 6141] = -'sd62923;
    data[ 6142] =  'sd51062;
    data[ 6143] =  'sd29752;
    data[ 6144] =  'sd44423;
    data[ 6145] = -'sd16721;
    data[ 6146] =  'sd46794;
    data[ 6147] = -'sd124;
    data[ 6148] = -'sd868;
    data[ 6149] = -'sd6076;
    data[ 6150] = -'sd42532;
    data[ 6151] =  'sd29958;
    data[ 6152] =  'sd45865;
    data[ 6153] = -'sd6627;
    data[ 6154] = -'sd46389;
    data[ 6155] =  'sd2959;
    data[ 6156] =  'sd20713;
    data[ 6157] = -'sd18850;
    data[ 6158] =  'sd31891;
    data[ 6159] =  'sd59396;
    data[ 6160] = -'sd75751;
    data[ 6161] = -'sd38734;
    data[ 6162] =  'sd56544;
    data[ 6163] =  'sd68126;
    data[ 6164] = -'sd14641;
    data[ 6165] =  'sd61354;
    data[ 6166] = -'sd62045;
    data[ 6167] =  'sd57208;
    data[ 6168] =  'sd72774;
    data[ 6169] =  'sd17895;
    data[ 6170] = -'sd38576;
    data[ 6171] =  'sd57650;
    data[ 6172] =  'sd75868;
    data[ 6173] =  'sd39553;
    data[ 6174] = -'sd50811;
    data[ 6175] = -'sd27995;
    data[ 6176] = -'sd32124;
    data[ 6177] = -'sd61027;
    data[ 6178] =  'sd64334;
    data[ 6179] = -'sd41185;
    data[ 6180] =  'sd39387;
    data[ 6181] = -'sd51973;
    data[ 6182] = -'sd36129;
    data[ 6183] =  'sd74779;
    data[ 6184] =  'sd31930;
    data[ 6185] =  'sd59669;
    data[ 6186] = -'sd73840;
    data[ 6187] = -'sd25357;
    data[ 6188] = -'sd13658;
    data[ 6189] =  'sd68235;
    data[ 6190] = -'sd13878;
    data[ 6191] =  'sd66695;
    data[ 6192] = -'sd24658;
    data[ 6193] = -'sd8765;
    data[ 6194] = -'sd61355;
    data[ 6195] =  'sd62038;
    data[ 6196] = -'sd57257;
    data[ 6197] = -'sd73117;
    data[ 6198] = -'sd20296;
    data[ 6199] =  'sd21769;
    data[ 6200] = -'sd11458;
    data[ 6201] = -'sd80206;
    data[ 6202] = -'sd69919;
    data[ 6203] =  'sd2090;
    data[ 6204] =  'sd14630;
    data[ 6205] = -'sd61431;
    data[ 6206] =  'sd61506;
    data[ 6207] = -'sd60981;
    data[ 6208] =  'sd64656;
    data[ 6209] = -'sd38931;
    data[ 6210] =  'sd55165;
    data[ 6211] =  'sd58473;
    data[ 6212] =  'sd81629;
    data[ 6213] =  'sd79880;
    data[ 6214] =  'sd67637;
    data[ 6215] = -'sd18064;
    data[ 6216] =  'sd37393;
    data[ 6217] = -'sd65931;
    data[ 6218] =  'sd30006;
    data[ 6219] =  'sd46201;
    data[ 6220] = -'sd4275;
    data[ 6221] = -'sd29925;
    data[ 6222] = -'sd45634;
    data[ 6223] =  'sd8244;
    data[ 6224] =  'sd57708;
    data[ 6225] =  'sd76274;
    data[ 6226] =  'sd42395;
    data[ 6227] = -'sd30917;
    data[ 6228] = -'sd52578;
    data[ 6229] = -'sd40364;
    data[ 6230] =  'sd45134;
    data[ 6231] = -'sd11744;
    data[ 6232] =  'sd81633;
    data[ 6233] =  'sd79908;
    data[ 6234] =  'sd67833;
    data[ 6235] = -'sd16692;
    data[ 6236] =  'sd46997;
    data[ 6237] =  'sd1297;
    data[ 6238] =  'sd9079;
    data[ 6239] =  'sd63553;
    data[ 6240] = -'sd46652;
    data[ 6241] =  'sd1118;
    data[ 6242] =  'sd7826;
    data[ 6243] =  'sd54782;
    data[ 6244] =  'sd55792;
    data[ 6245] =  'sd62862;
    data[ 6246] = -'sd51489;
    data[ 6247] = -'sd32741;
    data[ 6248] = -'sd65346;
    data[ 6249] =  'sd34101;
    data[ 6250] =  'sd74866;
    data[ 6251] =  'sd32539;
    data[ 6252] =  'sd63932;
    data[ 6253] = -'sd43999;
    data[ 6254] =  'sd19689;
    data[ 6255] = -'sd26018;
    data[ 6256] = -'sd18285;
    data[ 6257] =  'sd35846;
    data[ 6258] = -'sd76760;
    data[ 6259] = -'sd45797;
    data[ 6260] =  'sd7103;
    data[ 6261] =  'sd49721;
    data[ 6262] =  'sd20365;
    data[ 6263] = -'sd21286;
    data[ 6264] =  'sd14839;
    data[ 6265] = -'sd59968;
    data[ 6266] =  'sd71747;
    data[ 6267] =  'sd10706;
    data[ 6268] =  'sd74942;
    data[ 6269] =  'sd33071;
    data[ 6270] =  'sd67656;
    data[ 6271] = -'sd17931;
    data[ 6272] =  'sd38324;
    data[ 6273] = -'sd59414;
    data[ 6274] =  'sd75625;
    data[ 6275] =  'sd37852;
    data[ 6276] = -'sd62718;
    data[ 6277] =  'sd52497;
    data[ 6278] =  'sd39797;
    data[ 6279] = -'sd49103;
    data[ 6280] = -'sd16039;
    data[ 6281] =  'sd51568;
    data[ 6282] =  'sd33294;
    data[ 6283] =  'sd69217;
    data[ 6284] = -'sd7004;
    data[ 6285] = -'sd49028;
    data[ 6286] = -'sd15514;
    data[ 6287] =  'sd55243;
    data[ 6288] =  'sd59019;
    data[ 6289] = -'sd78390;
    data[ 6290] = -'sd57207;
    data[ 6291] = -'sd72767;
    data[ 6292] = -'sd17846;
    data[ 6293] =  'sd38919;
    data[ 6294] = -'sd55249;
    data[ 6295] = -'sd59061;
    data[ 6296] =  'sd78096;
    data[ 6297] =  'sd55149;
    data[ 6298] =  'sd58361;
    data[ 6299] =  'sd80845;
    data[ 6300] =  'sd74392;
    data[ 6301] =  'sd29221;
    data[ 6302] =  'sd40706;
    data[ 6303] = -'sd42740;
    data[ 6304] =  'sd28502;
    data[ 6305] =  'sd35673;
    data[ 6306] = -'sd77971;
    data[ 6307] = -'sd54274;
    data[ 6308] = -'sd52236;
    data[ 6309] = -'sd37970;
    data[ 6310] =  'sd61892;
    data[ 6311] = -'sd58279;
    data[ 6312] = -'sd80271;
    data[ 6313] = -'sd70374;
    data[ 6314] = -'sd1095;
    data[ 6315] = -'sd7665;
    data[ 6316] = -'sd53655;
    data[ 6317] = -'sd47903;
    data[ 6318] = -'sd7639;
    data[ 6319] = -'sd53473;
    data[ 6320] = -'sd46629;
    data[ 6321] =  'sd1279;
    data[ 6322] =  'sd8953;
    data[ 6323] =  'sd62671;
    data[ 6324] = -'sd52826;
    data[ 6325] = -'sd42100;
    data[ 6326] =  'sd32982;
    data[ 6327] =  'sd67033;
    data[ 6328] = -'sd22292;
    data[ 6329] =  'sd7797;
    data[ 6330] =  'sd54579;
    data[ 6331] =  'sd54371;
    data[ 6332] =  'sd52915;
    data[ 6333] =  'sd42723;
    data[ 6334] = -'sd28621;
    data[ 6335] = -'sd36506;
    data[ 6336] =  'sd72140;
    data[ 6337] =  'sd13457;
    data[ 6338] = -'sd69642;
    data[ 6339] =  'sd4029;
    data[ 6340] =  'sd28203;
    data[ 6341] =  'sd33580;
    data[ 6342] =  'sd71219;
    data[ 6343] =  'sd7010;
    data[ 6344] =  'sd49070;
    data[ 6345] =  'sd15808;
    data[ 6346] = -'sd53185;
    data[ 6347] = -'sd44613;
    data[ 6348] =  'sd15391;
    data[ 6349] = -'sd56104;
    data[ 6350] = -'sd65046;
    data[ 6351] =  'sd36201;
    data[ 6352] = -'sd74275;
    data[ 6353] = -'sd28402;
    data[ 6354] = -'sd34973;
    data[ 6355] = -'sd80970;
    data[ 6356] = -'sd75267;
    data[ 6357] = -'sd35346;
    data[ 6358] =  'sd80260;
    data[ 6359] =  'sd70297;
    data[ 6360] =  'sd556;
    data[ 6361] =  'sd3892;
    data[ 6362] =  'sd27244;
    data[ 6363] =  'sd26867;
    data[ 6364] =  'sd24228;
    data[ 6365] =  'sd5755;
    data[ 6366] =  'sd40285;
    data[ 6367] = -'sd45687;
    data[ 6368] =  'sd7873;
    data[ 6369] =  'sd55111;
    data[ 6370] =  'sd58095;
    data[ 6371] =  'sd78983;
    data[ 6372] =  'sd61358;
    data[ 6373] = -'sd62017;
    data[ 6374] =  'sd57404;
    data[ 6375] =  'sd74146;
    data[ 6376] =  'sd27499;
    data[ 6377] =  'sd28652;
    data[ 6378] =  'sd36723;
    data[ 6379] = -'sd70621;
    data[ 6380] = -'sd2824;
    data[ 6381] = -'sd19768;
    data[ 6382] =  'sd25465;
    data[ 6383] =  'sd14414;
    data[ 6384] = -'sd62943;
    data[ 6385] =  'sd50922;
    data[ 6386] =  'sd28772;
    data[ 6387] =  'sd37563;
    data[ 6388] = -'sd64741;
    data[ 6389] =  'sd38336;
    data[ 6390] = -'sd59330;
    data[ 6391] =  'sd76213;
    data[ 6392] =  'sd41968;
    data[ 6393] = -'sd33906;
    data[ 6394] = -'sd73501;
    data[ 6395] = -'sd22984;
    data[ 6396] =  'sd2953;
    data[ 6397] =  'sd20671;
    data[ 6398] = -'sd19144;
    data[ 6399] =  'sd29833;
    data[ 6400] =  'sd44990;
    data[ 6401] = -'sd12752;
    data[ 6402] =  'sd74577;
    data[ 6403] =  'sd30516;
    data[ 6404] =  'sd49771;
    data[ 6405] =  'sd20715;
    data[ 6406] = -'sd18836;
    data[ 6407] =  'sd31989;
    data[ 6408] =  'sd60082;
    data[ 6409] = -'sd70949;
    data[ 6410] = -'sd5120;
    data[ 6411] = -'sd35840;
    data[ 6412] =  'sd76802;
    data[ 6413] =  'sd46091;
    data[ 6414] = -'sd5045;
    data[ 6415] = -'sd35315;
    data[ 6416] =  'sd80477;
    data[ 6417] =  'sd71816;
    data[ 6418] =  'sd11189;
    data[ 6419] =  'sd78323;
    data[ 6420] =  'sd56738;
    data[ 6421] =  'sd69484;
    data[ 6422] = -'sd5135;
    data[ 6423] = -'sd35945;
    data[ 6424] =  'sd76067;
    data[ 6425] =  'sd40946;
    data[ 6426] = -'sd41060;
    data[ 6427] =  'sd40262;
    data[ 6428] = -'sd45848;
    data[ 6429] =  'sd6746;
    data[ 6430] =  'sd47222;
    data[ 6431] =  'sd2872;
    data[ 6432] =  'sd20104;
    data[ 6433] = -'sd23113;
    data[ 6434] =  'sd2050;
    data[ 6435] =  'sd14350;
    data[ 6436] = -'sd63391;
    data[ 6437] =  'sd47786;
    data[ 6438] =  'sd6820;
    data[ 6439] =  'sd47740;
    data[ 6440] =  'sd6498;
    data[ 6441] =  'sd45486;
    data[ 6442] = -'sd9280;
    data[ 6443] = -'sd64960;
    data[ 6444] =  'sd36803;
    data[ 6445] = -'sd70061;
    data[ 6446] =  'sd1096;
    data[ 6447] =  'sd7672;
    data[ 6448] =  'sd53704;
    data[ 6449] =  'sd48246;
    data[ 6450] =  'sd10040;
    data[ 6451] =  'sd70280;
    data[ 6452] =  'sd437;
    data[ 6453] =  'sd3059;
    data[ 6454] =  'sd21413;
    data[ 6455] = -'sd13950;
    data[ 6456] =  'sd66191;
    data[ 6457] = -'sd28186;
    data[ 6458] = -'sd33461;
    data[ 6459] = -'sd70386;
    data[ 6460] = -'sd1179;
    data[ 6461] = -'sd8253;
    data[ 6462] = -'sd57771;
    data[ 6463] = -'sd76715;
    data[ 6464] = -'sd45482;
    data[ 6465] =  'sd9308;
    data[ 6466] =  'sd65156;
    data[ 6467] = -'sd35431;
    data[ 6468] =  'sd79665;
    data[ 6469] =  'sd66132;
    data[ 6470] = -'sd28599;
    data[ 6471] = -'sd36352;
    data[ 6472] =  'sd73218;
    data[ 6473] =  'sd21003;
    data[ 6474] = -'sd16820;
    data[ 6475] =  'sd46101;
    data[ 6476] = -'sd4975;
    data[ 6477] = -'sd34825;
    data[ 6478] = -'sd79934;
    data[ 6479] = -'sd68015;
    data[ 6480] =  'sd15418;
    data[ 6481] = -'sd55915;
    data[ 6482] = -'sd63723;
    data[ 6483] =  'sd45462;
    data[ 6484] = -'sd9448;
    data[ 6485] = -'sd66136;
    data[ 6486] =  'sd28571;
    data[ 6487] =  'sd36156;
    data[ 6488] = -'sd74590;
    data[ 6489] = -'sd30607;
    data[ 6490] = -'sd50408;
    data[ 6491] = -'sd25174;
    data[ 6492] = -'sd12377;
    data[ 6493] =  'sd77202;
    data[ 6494] =  'sd48891;
    data[ 6495] =  'sd14555;
    data[ 6496] = -'sd61956;
    data[ 6497] =  'sd57831;
    data[ 6498] =  'sd77135;
    data[ 6499] =  'sd48422;
    data[ 6500] =  'sd11272;
    data[ 6501] =  'sd78904;
    data[ 6502] =  'sd60805;
    data[ 6503] = -'sd65888;
    data[ 6504] =  'sd30307;
    data[ 6505] =  'sd48308;
    data[ 6506] =  'sd10474;
    data[ 6507] =  'sd73318;
    data[ 6508] =  'sd21703;
    data[ 6509] = -'sd11920;
    data[ 6510] =  'sd80401;
    data[ 6511] =  'sd71284;
    data[ 6512] =  'sd7465;
    data[ 6513] =  'sd52255;
    data[ 6514] =  'sd38103;
    data[ 6515] = -'sd60961;
    data[ 6516] =  'sd64796;
    data[ 6517] = -'sd37951;
    data[ 6518] =  'sd62025;
    data[ 6519] = -'sd57348;
    data[ 6520] = -'sd73754;
    data[ 6521] = -'sd24755;
    data[ 6522] = -'sd9444;
    data[ 6523] = -'sd66108;
    data[ 6524] =  'sd28767;
    data[ 6525] =  'sd37528;
    data[ 6526] = -'sd64986;
    data[ 6527] =  'sd36621;
    data[ 6528] = -'sd71335;
    data[ 6529] = -'sd7822;
    data[ 6530] = -'sd54754;
    data[ 6531] = -'sd55596;
    data[ 6532] = -'sd61490;
    data[ 6533] =  'sd61093;
    data[ 6534] = -'sd63872;
    data[ 6535] =  'sd44419;
    data[ 6536] = -'sd16749;
    data[ 6537] =  'sd46598;
    data[ 6538] = -'sd1496;
    data[ 6539] = -'sd10472;
    data[ 6540] = -'sd73304;
    data[ 6541] = -'sd21605;
    data[ 6542] =  'sd12606;
    data[ 6543] = -'sd75599;
    data[ 6544] = -'sd37670;
    data[ 6545] =  'sd63992;
    data[ 6546] = -'sd43579;
    data[ 6547] =  'sd22629;
    data[ 6548] = -'sd5438;
    data[ 6549] = -'sd38066;
    data[ 6550] =  'sd61220;
    data[ 6551] = -'sd62983;
    data[ 6552] =  'sd50642;
    data[ 6553] =  'sd26812;
    data[ 6554] =  'sd23843;
    data[ 6555] =  'sd3060;
    data[ 6556] =  'sd21420;
    data[ 6557] = -'sd13901;
    data[ 6558] =  'sd66534;
    data[ 6559] = -'sd25785;
    data[ 6560] = -'sd16654;
    data[ 6561] =  'sd47263;
    data[ 6562] =  'sd3159;
    data[ 6563] =  'sd22113;
    data[ 6564] = -'sd9050;
    data[ 6565] = -'sd63350;
    data[ 6566] =  'sd48073;
    data[ 6567] =  'sd8829;
    data[ 6568] =  'sd61803;
    data[ 6569] = -'sd58902;
    data[ 6570] =  'sd79209;
    data[ 6571] =  'sd62940;
    data[ 6572] = -'sd50943;
    data[ 6573] = -'sd28919;
    data[ 6574] = -'sd38592;
    data[ 6575] =  'sd57538;
    data[ 6576] =  'sd75084;
    data[ 6577] =  'sd34065;
    data[ 6578] =  'sd74614;
    data[ 6579] =  'sd30775;
    data[ 6580] =  'sd51584;
    data[ 6581] =  'sd33406;
    data[ 6582] =  'sd70001;
    data[ 6583] = -'sd1516;
    data[ 6584] = -'sd10612;
    data[ 6585] = -'sd74284;
    data[ 6586] = -'sd28465;
    data[ 6587] = -'sd35414;
    data[ 6588] =  'sd79784;
    data[ 6589] =  'sd66965;
    data[ 6590] = -'sd22768;
    data[ 6591] =  'sd4465;
    data[ 6592] =  'sd31255;
    data[ 6593] =  'sd54944;
    data[ 6594] =  'sd56926;
    data[ 6595] =  'sd70800;
    data[ 6596] =  'sd4077;
    data[ 6597] =  'sd28539;
    data[ 6598] =  'sd35932;
    data[ 6599] = -'sd76158;
    data[ 6600] = -'sd41583;
    data[ 6601] =  'sd36601;
    data[ 6602] = -'sd71475;
    data[ 6603] = -'sd8802;
    data[ 6604] = -'sd61614;
    data[ 6605] =  'sd60225;
    data[ 6606] = -'sd69948;
    data[ 6607] =  'sd1887;
    data[ 6608] =  'sd13209;
    data[ 6609] = -'sd71378;
    data[ 6610] = -'sd8123;
    data[ 6611] = -'sd56861;
    data[ 6612] = -'sd70345;
    data[ 6613] = -'sd892;
    data[ 6614] = -'sd6244;
    data[ 6615] = -'sd43708;
    data[ 6616] =  'sd21726;
    data[ 6617] = -'sd11759;
    data[ 6618] =  'sd81528;
    data[ 6619] =  'sd79173;
    data[ 6620] =  'sd62688;
    data[ 6621] = -'sd52707;
    data[ 6622] = -'sd41267;
    data[ 6623] =  'sd38813;
    data[ 6624] = -'sd55991;
    data[ 6625] = -'sd64255;
    data[ 6626] =  'sd41738;
    data[ 6627] = -'sd35516;
    data[ 6628] =  'sd79070;
    data[ 6629] =  'sd61967;
    data[ 6630] = -'sd57754;
    data[ 6631] = -'sd76596;
    data[ 6632] = -'sd44649;
    data[ 6633] =  'sd15139;
    data[ 6634] = -'sd57868;
    data[ 6635] = -'sd77394;
    data[ 6636] = -'sd50235;
    data[ 6637] = -'sd23963;
    data[ 6638] = -'sd3900;
    data[ 6639] = -'sd27300;
    data[ 6640] = -'sd27259;
    data[ 6641] = -'sd26972;
    data[ 6642] = -'sd24963;
    data[ 6643] = -'sd10900;
    data[ 6644] = -'sd76300;
    data[ 6645] = -'sd42577;
    data[ 6646] =  'sd29643;
    data[ 6647] =  'sd43660;
    data[ 6648] = -'sd22062;
    data[ 6649] =  'sd9407;
    data[ 6650] =  'sd65849;
    data[ 6651] = -'sd30580;
    data[ 6652] = -'sd50219;
    data[ 6653] = -'sd23851;
    data[ 6654] = -'sd3116;
    data[ 6655] = -'sd21812;
    data[ 6656] =  'sd11157;
    data[ 6657] =  'sd78099;
    data[ 6658] =  'sd55170;
    data[ 6659] =  'sd58508;
    data[ 6660] =  'sd81874;
    data[ 6661] =  'sd81595;
    data[ 6662] =  'sd79642;
    data[ 6663] =  'sd65971;
    data[ 6664] = -'sd29726;
    data[ 6665] = -'sd44241;
    data[ 6666] =  'sd17995;
    data[ 6667] = -'sd37876;
    data[ 6668] =  'sd62550;
    data[ 6669] = -'sd53673;
    data[ 6670] = -'sd48029;
    data[ 6671] = -'sd8521;
    data[ 6672] = -'sd59647;
    data[ 6673] =  'sd73994;
    data[ 6674] =  'sd26435;
    data[ 6675] =  'sd21204;
    data[ 6676] = -'sd15413;
    data[ 6677] =  'sd55950;
    data[ 6678] =  'sd63968;
    data[ 6679] = -'sd43747;
    data[ 6680] =  'sd21453;
    data[ 6681] = -'sd13670;
    data[ 6682] =  'sd68151;
    data[ 6683] = -'sd14466;
    data[ 6684] =  'sd62579;
    data[ 6685] = -'sd53470;
    data[ 6686] = -'sd46608;
    data[ 6687] =  'sd1426;
    data[ 6688] =  'sd9982;
    data[ 6689] =  'sd69874;
    data[ 6690] = -'sd2405;
    data[ 6691] = -'sd16835;
    data[ 6692] =  'sd45996;
    data[ 6693] = -'sd5710;
    data[ 6694] = -'sd39970;
    data[ 6695] =  'sd47892;
    data[ 6696] =  'sd7562;
    data[ 6697] =  'sd52934;
    data[ 6698] =  'sd42856;
    data[ 6699] = -'sd27690;
    data[ 6700] = -'sd29989;
    data[ 6701] = -'sd46082;
    data[ 6702] =  'sd5108;
    data[ 6703] =  'sd35756;
    data[ 6704] = -'sd77390;
    data[ 6705] = -'sd50207;
    data[ 6706] = -'sd23767;
    data[ 6707] = -'sd2528;
    data[ 6708] = -'sd17696;
    data[ 6709] =  'sd39969;
    data[ 6710] = -'sd47899;
    data[ 6711] = -'sd7611;
    data[ 6712] = -'sd53277;
    data[ 6713] = -'sd45257;
    data[ 6714] =  'sd10883;
    data[ 6715] =  'sd76181;
    data[ 6716] =  'sd41744;
    data[ 6717] = -'sd35474;
    data[ 6718] =  'sd79364;
    data[ 6719] =  'sd64025;
    data[ 6720] = -'sd43348;
    data[ 6721] =  'sd24246;
    data[ 6722] =  'sd5881;
    data[ 6723] =  'sd41167;
    data[ 6724] = -'sd39513;
    data[ 6725] =  'sd51091;
    data[ 6726] =  'sd29955;
    data[ 6727] =  'sd45844;
    data[ 6728] = -'sd6774;
    data[ 6729] = -'sd47418;
    data[ 6730] = -'sd4244;
    data[ 6731] = -'sd29708;
    data[ 6732] = -'sd44115;
    data[ 6733] =  'sd18877;
    data[ 6734] = -'sd31702;
    data[ 6735] = -'sd58073;
    data[ 6736] = -'sd78829;
    data[ 6737] = -'sd60280;
    data[ 6738] =  'sd69563;
    data[ 6739] = -'sd4582;
    data[ 6740] = -'sd32074;
    data[ 6741] = -'sd60677;
    data[ 6742] =  'sd66784;
    data[ 6743] = -'sd24035;
    data[ 6744] = -'sd4404;
    data[ 6745] = -'sd30828;
    data[ 6746] = -'sd51955;
    data[ 6747] = -'sd36003;
    data[ 6748] =  'sd75661;
    data[ 6749] =  'sd38104;
    data[ 6750] = -'sd60954;
    data[ 6751] =  'sd64845;
    data[ 6752] = -'sd37608;
    data[ 6753] =  'sd64426;
    data[ 6754] = -'sd40541;
    data[ 6755] =  'sd43895;
    data[ 6756] = -'sd20417;
    data[ 6757] =  'sd20922;
    data[ 6758] = -'sd17387;
    data[ 6759] =  'sd42132;
    data[ 6760] = -'sd32758;
    data[ 6761] = -'sd65465;
    data[ 6762] =  'sd33268;
    data[ 6763] =  'sd69035;
    data[ 6764] = -'sd8278;
    data[ 6765] = -'sd57946;
    data[ 6766] = -'sd77940;
    data[ 6767] = -'sd54057;
    data[ 6768] = -'sd50717;
    data[ 6769] = -'sd27337;
    data[ 6770] = -'sd27518;
    data[ 6771] = -'sd28785;
    data[ 6772] = -'sd37654;
    data[ 6773] =  'sd64104;
    data[ 6774] = -'sd42795;
    data[ 6775] =  'sd28117;
    data[ 6776] =  'sd32978;
    data[ 6777] =  'sd67005;
    data[ 6778] = -'sd22488;
    data[ 6779] =  'sd6425;
    data[ 6780] =  'sd44975;
    data[ 6781] = -'sd12857;
    data[ 6782] =  'sd73842;
    data[ 6783] =  'sd25371;
    data[ 6784] =  'sd13756;
    data[ 6785] = -'sd67549;
    data[ 6786] =  'sd18680;
    data[ 6787] = -'sd33081;
    data[ 6788] = -'sd67726;
    data[ 6789] =  'sd17441;
    data[ 6790] = -'sd41754;
    data[ 6791] =  'sd35404;
    data[ 6792] = -'sd79854;
    data[ 6793] = -'sd67455;
    data[ 6794] =  'sd19338;
    data[ 6795] = -'sd28475;
    data[ 6796] = -'sd35484;
    data[ 6797] =  'sd79294;
    data[ 6798] =  'sd63535;
    data[ 6799] = -'sd46778;
    data[ 6800] =  'sd236;
    data[ 6801] =  'sd1652;
    data[ 6802] =  'sd11564;
    data[ 6803] =  'sd80948;
    data[ 6804] =  'sd75113;
    data[ 6805] =  'sd34268;
    data[ 6806] =  'sd76035;
    data[ 6807] =  'sd40722;
    data[ 6808] = -'sd42628;
    data[ 6809] =  'sd29286;
    data[ 6810] =  'sd41161;
    data[ 6811] = -'sd39555;
    data[ 6812] =  'sd50797;
    data[ 6813] =  'sd27897;
    data[ 6814] =  'sd31438;
    data[ 6815] =  'sd56225;
    data[ 6816] =  'sd65893;
    data[ 6817] = -'sd30272;
    data[ 6818] = -'sd48063;
    data[ 6819] = -'sd8759;
    data[ 6820] = -'sd61313;
    data[ 6821] =  'sd62332;
    data[ 6822] = -'sd55199;
    data[ 6823] = -'sd58711;
    data[ 6824] =  'sd80546;
    data[ 6825] =  'sd72299;
    data[ 6826] =  'sd14570;
    data[ 6827] = -'sd61851;
    data[ 6828] =  'sd58566;
    data[ 6829] = -'sd81561;
    data[ 6830] = -'sd79404;
    data[ 6831] = -'sd64305;
    data[ 6832] =  'sd41388;
    data[ 6833] = -'sd37966;
    data[ 6834] =  'sd61920;
    data[ 6835] = -'sd58083;
    data[ 6836] = -'sd78899;
    data[ 6837] = -'sd60770;
    data[ 6838] =  'sd66133;
    data[ 6839] = -'sd28592;
    data[ 6840] = -'sd36303;
    data[ 6841] =  'sd73561;
    data[ 6842] =  'sd23404;
    data[ 6843] = -'sd13;
    data[ 6844] = -'sd91;
    data[ 6845] = -'sd637;
    data[ 6846] = -'sd4459;
    data[ 6847] = -'sd31213;
    data[ 6848] = -'sd54650;
    data[ 6849] = -'sd54868;
    data[ 6850] = -'sd56394;
    data[ 6851] = -'sd67076;
    data[ 6852] =  'sd21991;
    data[ 6853] = -'sd9904;
    data[ 6854] = -'sd69328;
    data[ 6855] =  'sd6227;
    data[ 6856] =  'sd43589;
    data[ 6857] = -'sd22559;
    data[ 6858] =  'sd5928;
    data[ 6859] =  'sd41496;
    data[ 6860] = -'sd37210;
    data[ 6861] =  'sd67212;
    data[ 6862] = -'sd21039;
    data[ 6863] =  'sd16568;
    data[ 6864] = -'sd47865;
    data[ 6865] = -'sd7373;
    data[ 6866] = -'sd51611;
    data[ 6867] = -'sd33595;
    data[ 6868] = -'sd71324;
    data[ 6869] = -'sd7745;
    data[ 6870] = -'sd54215;
    data[ 6871] = -'sd51823;
    data[ 6872] = -'sd35079;
    data[ 6873] = -'sd81712;
    data[ 6874] = -'sd80461;
    data[ 6875] = -'sd71704;
    data[ 6876] = -'sd10405;
    data[ 6877] = -'sd72835;
    data[ 6878] = -'sd18322;
    data[ 6879] =  'sd35587;
    data[ 6880] = -'sd78573;
    data[ 6881] = -'sd58488;
    data[ 6882] = -'sd81734;
    data[ 6883] = -'sd80615;
    data[ 6884] = -'sd72782;
    data[ 6885] = -'sd17951;
    data[ 6886] =  'sd38184;
    data[ 6887] = -'sd60394;
    data[ 6888] =  'sd68765;
    data[ 6889] = -'sd10168;
    data[ 6890] = -'sd71176;
    data[ 6891] = -'sd6709;
    data[ 6892] = -'sd46963;
    data[ 6893] = -'sd1059;
    data[ 6894] = -'sd7413;
    data[ 6895] = -'sd51891;
    data[ 6896] = -'sd35555;
    data[ 6897] =  'sd78797;
    data[ 6898] =  'sd60056;
    data[ 6899] = -'sd71131;
    data[ 6900] = -'sd6394;
    data[ 6901] = -'sd44758;
    data[ 6902] =  'sd14376;
    data[ 6903] = -'sd63209;
    data[ 6904] =  'sd49060;
    data[ 6905] =  'sd15738;
    data[ 6906] = -'sd53675;
    data[ 6907] = -'sd48043;
    data[ 6908] = -'sd8619;
    data[ 6909] = -'sd60333;
    data[ 6910] =  'sd69192;
    data[ 6911] = -'sd7179;
    data[ 6912] = -'sd50253;
    data[ 6913] = -'sd24089;
    data[ 6914] = -'sd4782;
    data[ 6915] = -'sd33474;
    data[ 6916] = -'sd70477;
    data[ 6917] = -'sd1816;
    data[ 6918] = -'sd12712;
    data[ 6919] =  'sd74857;
    data[ 6920] =  'sd32476;
    data[ 6921] =  'sd63491;
    data[ 6922] = -'sd47086;
    data[ 6923] = -'sd1920;
    data[ 6924] = -'sd13440;
    data[ 6925] =  'sd69761;
    data[ 6926] = -'sd3196;
    data[ 6927] = -'sd22372;
    data[ 6928] =  'sd7237;
    data[ 6929] =  'sd50659;
    data[ 6930] =  'sd26931;
    data[ 6931] =  'sd24676;
    data[ 6932] =  'sd8891;
    data[ 6933] =  'sd62237;
    data[ 6934] = -'sd55864;
    data[ 6935] = -'sd63366;
    data[ 6936] =  'sd47961;
    data[ 6937] =  'sd8045;
    data[ 6938] =  'sd56315;
    data[ 6939] =  'sd66523;
    data[ 6940] = -'sd25862;
    data[ 6941] = -'sd17193;
    data[ 6942] =  'sd43490;
    data[ 6943] = -'sd23252;
    data[ 6944] =  'sd1077;
    data[ 6945] =  'sd7539;
    data[ 6946] =  'sd52773;
    data[ 6947] =  'sd41729;
    data[ 6948] = -'sd35579;
    data[ 6949] =  'sd78629;
    data[ 6950] =  'sd58880;
    data[ 6951] = -'sd79363;
    data[ 6952] = -'sd64018;
    data[ 6953] =  'sd43397;
    data[ 6954] = -'sd23903;
    data[ 6955] = -'sd3480;
    data[ 6956] = -'sd24360;
    data[ 6957] = -'sd6679;
    data[ 6958] = -'sd46753;
    data[ 6959] =  'sd411;
    data[ 6960] =  'sd2877;
    data[ 6961] =  'sd20139;
    data[ 6962] = -'sd22868;
    data[ 6963] =  'sd3765;
    data[ 6964] =  'sd26355;
    data[ 6965] =  'sd20644;
    data[ 6966] = -'sd19333;
    data[ 6967] =  'sd28510;
    data[ 6968] =  'sd35729;
    data[ 6969] = -'sd77579;
    data[ 6970] = -'sd51530;
    data[ 6971] = -'sd33028;
    data[ 6972] = -'sd67355;
    data[ 6973] =  'sd20038;
    data[ 6974] = -'sd23575;
    data[ 6975] = -'sd1184;
    data[ 6976] = -'sd8288;
    data[ 6977] = -'sd58016;
    data[ 6978] = -'sd78430;
    data[ 6979] = -'sd57487;
    data[ 6980] = -'sd74727;
    data[ 6981] = -'sd31566;
    data[ 6982] = -'sd57121;
    data[ 6983] = -'sd72165;
    data[ 6984] = -'sd13632;
    data[ 6985] =  'sd68417;
    data[ 6986] = -'sd12604;
    data[ 6987] =  'sd75613;
    data[ 6988] =  'sd37768;
    data[ 6989] = -'sd63306;
    data[ 6990] =  'sd48381;
    data[ 6991] =  'sd10985;
    data[ 6992] =  'sd76895;
    data[ 6993] =  'sd46742;
    data[ 6994] = -'sd488;
    data[ 6995] = -'sd3416;
    data[ 6996] = -'sd23912;
    data[ 6997] = -'sd3543;
    data[ 6998] = -'sd24801;
    data[ 6999] = -'sd9766;
    data[ 7000] = -'sd68362;
    data[ 7001] =  'sd12989;
    data[ 7002] = -'sd72918;
    data[ 7003] = -'sd18903;
    data[ 7004] =  'sd31520;
    data[ 7005] =  'sd56799;
    data[ 7006] =  'sd69911;
    data[ 7007] = -'sd2146;
    data[ 7008] = -'sd15022;
    data[ 7009] =  'sd58687;
    data[ 7010] = -'sd80714;
    data[ 7011] = -'sd73475;
    data[ 7012] = -'sd22802;
    data[ 7013] =  'sd4227;
    data[ 7014] =  'sd29589;
    data[ 7015] =  'sd43282;
    data[ 7016] = -'sd24708;
    data[ 7017] = -'sd9115;
    data[ 7018] = -'sd63805;
    data[ 7019] =  'sd44888;
    data[ 7020] = -'sd13466;
    data[ 7021] =  'sd69579;
    data[ 7022] = -'sd4470;
    data[ 7023] = -'sd31290;
    data[ 7024] = -'sd55189;
    data[ 7025] = -'sd58641;
    data[ 7026] =  'sd81036;
    data[ 7027] =  'sd75729;
    data[ 7028] =  'sd38580;
    data[ 7029] = -'sd57622;
    data[ 7030] = -'sd75672;
    data[ 7031] = -'sd38181;
    data[ 7032] =  'sd60415;
    data[ 7033] = -'sd68618;
    data[ 7034] =  'sd11197;
    data[ 7035] =  'sd78379;
    data[ 7036] =  'sd57130;
    data[ 7037] =  'sd72228;
    data[ 7038] =  'sd14073;
    data[ 7039] = -'sd65330;
    data[ 7040] =  'sd34213;
    data[ 7041] =  'sd75650;
    data[ 7042] =  'sd38027;
    data[ 7043] = -'sd61493;
    data[ 7044] =  'sd61072;
    data[ 7045] = -'sd64019;
    data[ 7046] =  'sd43390;
    data[ 7047] = -'sd23952;
    data[ 7048] = -'sd3823;
    data[ 7049] = -'sd26761;
    data[ 7050] = -'sd23486;
    data[ 7051] = -'sd561;
    data[ 7052] = -'sd3927;
    data[ 7053] = -'sd27489;
    data[ 7054] = -'sd28582;
    data[ 7055] = -'sd36233;
    data[ 7056] =  'sd74051;
    data[ 7057] =  'sd26834;
    data[ 7058] =  'sd23997;
    data[ 7059] =  'sd4138;
    data[ 7060] =  'sd28966;
    data[ 7061] =  'sd38921;
    data[ 7062] = -'sd55235;
    data[ 7063] = -'sd58963;
    data[ 7064] =  'sd78782;
    data[ 7065] =  'sd59951;
    data[ 7066] = -'sd71866;
    data[ 7067] = -'sd11539;
    data[ 7068] = -'sd80773;
    data[ 7069] = -'sd73888;
    data[ 7070] = -'sd25693;
    data[ 7071] = -'sd16010;
    data[ 7072] =  'sd51771;
    data[ 7073] =  'sd34715;
    data[ 7074] =  'sd79164;
    data[ 7075] =  'sd62625;
    data[ 7076] = -'sd53148;
    data[ 7077] = -'sd44354;
    data[ 7078] =  'sd17204;
    data[ 7079] = -'sd43413;
    data[ 7080] =  'sd23791;
    data[ 7081] =  'sd2696;
    data[ 7082] =  'sd18872;
    data[ 7083] = -'sd31737;
    data[ 7084] = -'sd58318;
    data[ 7085] = -'sd80544;
    data[ 7086] = -'sd72285;
    data[ 7087] = -'sd14472;
    data[ 7088] =  'sd62537;
    data[ 7089] = -'sd53764;
    data[ 7090] = -'sd48666;
    data[ 7091] = -'sd12980;
    data[ 7092] =  'sd72981;
    data[ 7093] =  'sd19344;
    data[ 7094] = -'sd28433;
    data[ 7095] = -'sd35190;
    data[ 7096] =  'sd81352;
    data[ 7097] =  'sd77941;
    data[ 7098] =  'sd54064;
    data[ 7099] =  'sd50766;
    data[ 7100] =  'sd27680;
    data[ 7101] =  'sd29919;
    data[ 7102] =  'sd45592;
    data[ 7103] = -'sd8538;
    data[ 7104] = -'sd59766;
    data[ 7105] =  'sd73161;
    data[ 7106] =  'sd20604;
    data[ 7107] = -'sd19613;
    data[ 7108] =  'sd26550;
    data[ 7109] =  'sd22009;
    data[ 7110] = -'sd9778;
    data[ 7111] = -'sd68446;
    data[ 7112] =  'sd12401;
    data[ 7113] = -'sd77034;
    data[ 7114] = -'sd47715;
    data[ 7115] = -'sd6323;
    data[ 7116] = -'sd44261;
    data[ 7117] =  'sd17855;
    data[ 7118] = -'sd38856;
    data[ 7119] =  'sd55690;
    data[ 7120] =  'sd62148;
    data[ 7121] = -'sd56487;
    data[ 7122] = -'sd67727;
    data[ 7123] =  'sd17434;
    data[ 7124] = -'sd41803;
    data[ 7125] =  'sd35061;
    data[ 7126] =  'sd81586;
    data[ 7127] =  'sd79579;
    data[ 7128] =  'sd65530;
    data[ 7129] = -'sd32813;
    data[ 7130] = -'sd65850;
    data[ 7131] =  'sd30573;
    data[ 7132] =  'sd50170;
    data[ 7133] =  'sd23508;
    data[ 7134] =  'sd715;
    data[ 7135] =  'sd5005;
    data[ 7136] =  'sd35035;
    data[ 7137] =  'sd81404;
    data[ 7138] =  'sd78305;
    data[ 7139] =  'sd56612;
    data[ 7140] =  'sd68602;
    data[ 7141] = -'sd11309;
    data[ 7142] = -'sd79163;
    data[ 7143] = -'sd62618;
    data[ 7144] =  'sd53197;
    data[ 7145] =  'sd44697;
    data[ 7146] = -'sd14803;
    data[ 7147] =  'sd60220;
    data[ 7148] = -'sd69983;
    data[ 7149] =  'sd1642;
    data[ 7150] =  'sd11494;
    data[ 7151] =  'sd80458;
    data[ 7152] =  'sd71683;
    data[ 7153] =  'sd10258;
    data[ 7154] =  'sd71806;
    data[ 7155] =  'sd11119;
    data[ 7156] =  'sd77833;
    data[ 7157] =  'sd53308;
    data[ 7158] =  'sd45474;
    data[ 7159] = -'sd9364;
    data[ 7160] = -'sd65548;
    data[ 7161] =  'sd32687;
    data[ 7162] =  'sd64968;
    data[ 7163] = -'sd36747;
    data[ 7164] =  'sd70453;
    data[ 7165] =  'sd1648;
    data[ 7166] =  'sd11536;
    data[ 7167] =  'sd80752;
    data[ 7168] =  'sd73741;
    data[ 7169] =  'sd24664;
    data[ 7170] =  'sd8807;
    data[ 7171] =  'sd61649;
    data[ 7172] = -'sd59980;
    data[ 7173] =  'sd71663;
    data[ 7174] =  'sd10118;
    data[ 7175] =  'sd70826;
    data[ 7176] =  'sd4259;
    data[ 7177] =  'sd29813;
    data[ 7178] =  'sd44850;
    data[ 7179] = -'sd13732;
    data[ 7180] =  'sd67717;
    data[ 7181] = -'sd17504;
    data[ 7182] =  'sd41313;
    data[ 7183] = -'sd38491;
    data[ 7184] =  'sd58245;
    data[ 7185] =  'sd80033;
    data[ 7186] =  'sd68708;
    data[ 7187] = -'sd10567;
    data[ 7188] = -'sd73969;
    data[ 7189] = -'sd26260;
    data[ 7190] = -'sd19979;
    data[ 7191] =  'sd23988;
    data[ 7192] =  'sd4075;
    data[ 7193] =  'sd28525;
    data[ 7194] =  'sd35834;
    data[ 7195] = -'sd76844;
    data[ 7196] = -'sd46385;
    data[ 7197] =  'sd2987;
    data[ 7198] =  'sd20909;
    data[ 7199] = -'sd17478;
    data[ 7200] =  'sd41495;
    data[ 7201] = -'sd37217;
    data[ 7202] =  'sd67163;
    data[ 7203] = -'sd21382;
    data[ 7204] =  'sd14167;
    data[ 7205] = -'sd64672;
    data[ 7206] =  'sd38819;
    data[ 7207] = -'sd55949;
    data[ 7208] = -'sd63961;
    data[ 7209] =  'sd43796;
    data[ 7210] = -'sd21110;
    data[ 7211] =  'sd16071;
    data[ 7212] = -'sd51344;
    data[ 7213] = -'sd31726;
    data[ 7214] = -'sd58241;
    data[ 7215] = -'sd80005;
    data[ 7216] = -'sd68512;
    data[ 7217] =  'sd11939;
    data[ 7218] = -'sd80268;
    data[ 7219] = -'sd70353;
    data[ 7220] = -'sd948;
    data[ 7221] = -'sd6636;
    data[ 7222] = -'sd46452;
    data[ 7223] =  'sd2518;
    data[ 7224] =  'sd17626;
    data[ 7225] = -'sd40459;
    data[ 7226] =  'sd44469;
    data[ 7227] = -'sd16399;
    data[ 7228] =  'sd49048;
    data[ 7229] =  'sd15654;
    data[ 7230] = -'sd54263;
    data[ 7231] = -'sd52159;
    data[ 7232] = -'sd37431;
    data[ 7233] =  'sd65665;
    data[ 7234] = -'sd31868;
    data[ 7235] = -'sd59235;
    data[ 7236] =  'sd76878;
    data[ 7237] =  'sd46623;
    data[ 7238] = -'sd1321;
    data[ 7239] = -'sd9247;
    data[ 7240] = -'sd64729;
    data[ 7241] =  'sd38420;
    data[ 7242] = -'sd58742;
    data[ 7243] =  'sd80329;
    data[ 7244] =  'sd70780;
    data[ 7245] =  'sd3937;
    data[ 7246] =  'sd27559;
    data[ 7247] =  'sd29072;
    data[ 7248] =  'sd39663;
    data[ 7249] = -'sd50041;
    data[ 7250] = -'sd22605;
    data[ 7251] =  'sd5606;
    data[ 7252] =  'sd39242;
    data[ 7253] = -'sd52988;
    data[ 7254] = -'sd43234;
    data[ 7255] =  'sd25044;
    data[ 7256] =  'sd11467;
    data[ 7257] =  'sd80269;
    data[ 7258] =  'sd70360;
    data[ 7259] =  'sd997;
    data[ 7260] =  'sd6979;
    data[ 7261] =  'sd48853;
    data[ 7262] =  'sd14289;
    data[ 7263] = -'sd63818;
    data[ 7264] =  'sd44797;
    data[ 7265] = -'sd14103;
    data[ 7266] =  'sd65120;
    data[ 7267] = -'sd35683;
    data[ 7268] =  'sd77901;
    data[ 7269] =  'sd53784;
    data[ 7270] =  'sd48806;
    data[ 7271] =  'sd13960;
    data[ 7272] = -'sd66121;
    data[ 7273] =  'sd28676;
    data[ 7274] =  'sd36891;
    data[ 7275] = -'sd69445;
    data[ 7276] =  'sd5408;
    data[ 7277] =  'sd37856;
    data[ 7278] = -'sd62690;
    data[ 7279] =  'sd52693;
    data[ 7280] =  'sd41169;
    data[ 7281] = -'sd39499;
    data[ 7282] =  'sd51189;
    data[ 7283] =  'sd30641;
    data[ 7284] =  'sd50646;
    data[ 7285] =  'sd26840;
    data[ 7286] =  'sd24039;
    data[ 7287] =  'sd4432;
    data[ 7288] =  'sd31024;
    data[ 7289] =  'sd53327;
    data[ 7290] =  'sd45607;
    data[ 7291] = -'sd8433;
    data[ 7292] = -'sd59031;
    data[ 7293] =  'sd78306;
    data[ 7294] =  'sd56619;
    data[ 7295] =  'sd68651;
    data[ 7296] = -'sd10966;
    data[ 7297] = -'sd76762;
    data[ 7298] = -'sd45811;
    data[ 7299] =  'sd7005;
    data[ 7300] =  'sd49035;
    data[ 7301] =  'sd15563;
    data[ 7302] = -'sd54900;
    data[ 7303] = -'sd56618;
    data[ 7304] = -'sd68644;
    data[ 7305] =  'sd11015;
    data[ 7306] =  'sd77105;
    data[ 7307] =  'sd48212;
    data[ 7308] =  'sd9802;
    data[ 7309] =  'sd68614;
    data[ 7310] = -'sd11225;
    data[ 7311] = -'sd78575;
    data[ 7312] = -'sd58502;
    data[ 7313] = -'sd81832;
    data[ 7314] = -'sd81301;
    data[ 7315] = -'sd77584;
    data[ 7316] = -'sd51565;
    data[ 7317] = -'sd33273;
    data[ 7318] = -'sd69070;
    data[ 7319] =  'sd8033;
    data[ 7320] =  'sd56231;
    data[ 7321] =  'sd65935;
    data[ 7322] = -'sd29978;
    data[ 7323] = -'sd46005;
    data[ 7324] =  'sd5647;
    data[ 7325] =  'sd39529;
    data[ 7326] = -'sd50979;
    data[ 7327] = -'sd29171;
    data[ 7328] = -'sd40356;
    data[ 7329] =  'sd45190;
    data[ 7330] = -'sd11352;
    data[ 7331] = -'sd79464;
    data[ 7332] = -'sd64725;
    data[ 7333] =  'sd38448;
    data[ 7334] = -'sd58546;
    data[ 7335] =  'sd81701;
    data[ 7336] =  'sd80384;
    data[ 7337] =  'sd71165;
    data[ 7338] =  'sd6632;
    data[ 7339] =  'sd46424;
    data[ 7340] = -'sd2714;
    data[ 7341] = -'sd18998;
    data[ 7342] =  'sd30855;
    data[ 7343] =  'sd52144;
    data[ 7344] =  'sd37326;
    data[ 7345] = -'sd66400;
    data[ 7346] =  'sd26723;
    data[ 7347] =  'sd23220;
    data[ 7348] = -'sd1301;
    data[ 7349] = -'sd9107;
    data[ 7350] = -'sd63749;
    data[ 7351] =  'sd45280;
    data[ 7352] = -'sd10722;
    data[ 7353] = -'sd75054;
    data[ 7354] = -'sd33855;
    data[ 7355] = -'sd73144;
    data[ 7356] = -'sd20485;
    data[ 7357] =  'sd20446;
    data[ 7358] = -'sd20719;
    data[ 7359] =  'sd18808;
    data[ 7360] = -'sd32185;
    data[ 7361] = -'sd61454;
    data[ 7362] =  'sd61345;
    data[ 7363] = -'sd62108;
    data[ 7364] =  'sd56767;
    data[ 7365] =  'sd69687;
    data[ 7366] = -'sd3714;
    data[ 7367] = -'sd25998;
    data[ 7368] = -'sd18145;
    data[ 7369] =  'sd36826;
    data[ 7370] = -'sd69900;
    data[ 7371] =  'sd2223;
    data[ 7372] =  'sd15561;
    data[ 7373] = -'sd54914;
    data[ 7374] = -'sd56716;
    data[ 7375] = -'sd69330;
    data[ 7376] =  'sd6213;
    data[ 7377] =  'sd43491;
    data[ 7378] = -'sd23245;
    data[ 7379] =  'sd1126;
    data[ 7380] =  'sd7882;
    data[ 7381] =  'sd55174;
    data[ 7382] =  'sd58536;
    data[ 7383] = -'sd81771;
    data[ 7384] = -'sd80874;
    data[ 7385] = -'sd74595;
    data[ 7386] = -'sd30642;
    data[ 7387] = -'sd50653;
    data[ 7388] = -'sd26889;
    data[ 7389] = -'sd24382;
    data[ 7390] = -'sd6833;
    data[ 7391] = -'sd47831;
    data[ 7392] = -'sd7135;
    data[ 7393] = -'sd49945;
    data[ 7394] = -'sd21933;
    data[ 7395] =  'sd10310;
    data[ 7396] =  'sd72170;
    data[ 7397] =  'sd13667;
    data[ 7398] = -'sd68172;
    data[ 7399] =  'sd14319;
    data[ 7400] = -'sd63608;
    data[ 7401] =  'sd46267;
    data[ 7402] = -'sd3813;
    data[ 7403] = -'sd26691;
    data[ 7404] = -'sd22996;
    data[ 7405] =  'sd2869;
    data[ 7406] =  'sd20083;
    data[ 7407] = -'sd23260;
    data[ 7408] =  'sd1021;
    data[ 7409] =  'sd7147;
    data[ 7410] =  'sd50029;
    data[ 7411] =  'sd22521;
    data[ 7412] = -'sd6194;
    data[ 7413] = -'sd43358;
    data[ 7414] =  'sd24176;
    data[ 7415] =  'sd5391;
    data[ 7416] =  'sd37737;
    data[ 7417] = -'sd63523;
    data[ 7418] =  'sd46862;
    data[ 7419] =  'sd352;
    data[ 7420] =  'sd2464;
    data[ 7421] =  'sd17248;
    data[ 7422] = -'sd43105;
    data[ 7423] =  'sd25947;
    data[ 7424] =  'sd17788;
    data[ 7425] = -'sd39325;
    data[ 7426] =  'sd52407;
    data[ 7427] =  'sd39167;
    data[ 7428] = -'sd53513;
    data[ 7429] = -'sd46909;
    data[ 7430] = -'sd681;
    data[ 7431] = -'sd4767;
    data[ 7432] = -'sd33369;
    data[ 7433] = -'sd69742;
    data[ 7434] =  'sd3329;
    data[ 7435] =  'sd23303;
    data[ 7436] = -'sd720;
    data[ 7437] = -'sd5040;
    data[ 7438] = -'sd35280;
    data[ 7439] =  'sd80722;
    data[ 7440] =  'sd73531;
    data[ 7441] =  'sd23194;
    data[ 7442] = -'sd1483;
    data[ 7443] = -'sd10381;
    data[ 7444] = -'sd72667;
    data[ 7445] = -'sd17146;
    data[ 7446] =  'sd43819;
    data[ 7447] = -'sd20949;
    data[ 7448] =  'sd17198;
    data[ 7449] = -'sd43455;
    data[ 7450] =  'sd23497;
    data[ 7451] =  'sd638;
    data[ 7452] =  'sd4466;
    data[ 7453] =  'sd31262;
    data[ 7454] =  'sd54993;
    data[ 7455] =  'sd57269;
    data[ 7456] =  'sd73201;
    data[ 7457] =  'sd20884;
    data[ 7458] = -'sd17653;
    data[ 7459] =  'sd40270;
    data[ 7460] = -'sd45792;
    data[ 7461] =  'sd7138;
    data[ 7462] =  'sd49966;
    data[ 7463] =  'sd22080;
    data[ 7464] = -'sd9281;
    data[ 7465] = -'sd64967;
    data[ 7466] =  'sd36754;
    data[ 7467] = -'sd70404;
    data[ 7468] = -'sd1305;
    data[ 7469] = -'sd9135;
    data[ 7470] = -'sd63945;
    data[ 7471] =  'sd43908;
    data[ 7472] = -'sd20326;
    data[ 7473] =  'sd21559;
    data[ 7474] = -'sd12928;
    data[ 7475] =  'sd73345;
    data[ 7476] =  'sd21892;
    data[ 7477] = -'sd10597;
    data[ 7478] = -'sd74179;
    data[ 7479] = -'sd27730;
    data[ 7480] = -'sd30269;
    data[ 7481] = -'sd48042;
    data[ 7482] = -'sd8612;
    data[ 7483] = -'sd60284;
    data[ 7484] =  'sd69535;
    data[ 7485] = -'sd4778;
    data[ 7486] = -'sd33446;
    data[ 7487] = -'sd70281;
    data[ 7488] = -'sd444;
    data[ 7489] = -'sd3108;
    data[ 7490] = -'sd21756;
    data[ 7491] =  'sd11549;
    data[ 7492] =  'sd80843;
    data[ 7493] =  'sd74378;
    data[ 7494] =  'sd29123;
    data[ 7495] =  'sd40020;
    data[ 7496] = -'sd47542;
    data[ 7497] = -'sd5112;
    data[ 7498] = -'sd35784;
    data[ 7499] =  'sd77194;
    data[ 7500] =  'sd48835;
    data[ 7501] =  'sd14163;
    data[ 7502] = -'sd64700;
    data[ 7503] =  'sd38623;
    data[ 7504] = -'sd57321;
    data[ 7505] = -'sd73565;
    data[ 7506] = -'sd23432;
    data[ 7507] = -'sd183;
    data[ 7508] = -'sd1281;
    data[ 7509] = -'sd8967;
    data[ 7510] = -'sd62769;
    data[ 7511] =  'sd52140;
    data[ 7512] =  'sd37298;
    data[ 7513] = -'sd66596;
    data[ 7514] =  'sd25351;
    data[ 7515] =  'sd13616;
    data[ 7516] = -'sd68529;
    data[ 7517] =  'sd11820;
    data[ 7518] = -'sd81101;
    data[ 7519] = -'sd76184;
    data[ 7520] = -'sd41765;
    data[ 7521] =  'sd35327;
    data[ 7522] = -'sd80393;
    data[ 7523] = -'sd71228;
    data[ 7524] = -'sd7073;
    data[ 7525] = -'sd49511;
    data[ 7526] = -'sd18895;
    data[ 7527] =  'sd31576;
    data[ 7528] =  'sd57191;
    data[ 7529] =  'sd72655;
    data[ 7530] =  'sd17062;
    data[ 7531] = -'sd44407;
    data[ 7532] =  'sd16833;
    data[ 7533] = -'sd46010;
    data[ 7534] =  'sd5612;
    data[ 7535] =  'sd39284;
    data[ 7536] = -'sd52694;
    data[ 7537] = -'sd41176;
    data[ 7538] =  'sd39450;
    data[ 7539] = -'sd51532;
    data[ 7540] = -'sd33042;
    data[ 7541] = -'sd67453;
    data[ 7542] =  'sd19352;
    data[ 7543] = -'sd28377;
    data[ 7544] = -'sd34798;
    data[ 7545] = -'sd79745;
    data[ 7546] = -'sd66692;
    data[ 7547] =  'sd24679;
    data[ 7548] =  'sd8912;
    data[ 7549] =  'sd62384;
    data[ 7550] = -'sd54835;
    data[ 7551] = -'sd56163;
    data[ 7552] = -'sd65459;
    data[ 7553] =  'sd33310;
    data[ 7554] =  'sd69329;
    data[ 7555] = -'sd6220;
    data[ 7556] = -'sd43540;
    data[ 7557] =  'sd22902;
    data[ 7558] = -'sd3527;
    data[ 7559] = -'sd24689;
    data[ 7560] = -'sd8982;
    data[ 7561] = -'sd62874;
    data[ 7562] =  'sd51405;
    data[ 7563] =  'sd32153;
    data[ 7564] =  'sd61230;
    data[ 7565] = -'sd62913;
    data[ 7566] =  'sd51132;
    data[ 7567] =  'sd30242;
    data[ 7568] =  'sd47853;
    data[ 7569] =  'sd7289;
    data[ 7570] =  'sd51023;
    data[ 7571] =  'sd29479;
    data[ 7572] =  'sd42512;
    data[ 7573] = -'sd30098;
    data[ 7574] = -'sd46845;
    data[ 7575] = -'sd233;
    data[ 7576] = -'sd1631;
    data[ 7577] = -'sd11417;
    data[ 7578] = -'sd79919;
    data[ 7579] = -'sd67910;
    data[ 7580] =  'sd16153;
    data[ 7581] = -'sd50770;
    data[ 7582] = -'sd27708;
    data[ 7583] = -'sd30115;
    data[ 7584] = -'sd46964;
    data[ 7585] = -'sd1066;
    data[ 7586] = -'sd7462;
    data[ 7587] = -'sd52234;
    data[ 7588] = -'sd37956;
    data[ 7589] =  'sd61990;
    data[ 7590] = -'sd57593;
    data[ 7591] = -'sd75469;
    data[ 7592] = -'sd36760;
    data[ 7593] =  'sd70362;
    data[ 7594] =  'sd1011;
    data[ 7595] =  'sd7077;
    data[ 7596] =  'sd49539;
    data[ 7597] =  'sd19091;
    data[ 7598] = -'sd30204;
    data[ 7599] = -'sd47587;
    data[ 7600] = -'sd5427;
    data[ 7601] = -'sd37989;
    data[ 7602] =  'sd61759;
    data[ 7603] = -'sd59210;
    data[ 7604] =  'sd77053;
    data[ 7605] =  'sd47848;
    data[ 7606] =  'sd7254;
    data[ 7607] =  'sd50778;
    data[ 7608] =  'sd27764;
    data[ 7609] =  'sd30507;
    data[ 7610] =  'sd49708;
    data[ 7611] =  'sd20274;
    data[ 7612] = -'sd21923;
    data[ 7613] =  'sd10380;
    data[ 7614] =  'sd72660;
    data[ 7615] =  'sd17097;
    data[ 7616] = -'sd44162;
    data[ 7617] =  'sd18548;
    data[ 7618] = -'sd34005;
    data[ 7619] = -'sd74194;
    data[ 7620] = -'sd27835;
    data[ 7621] = -'sd31004;
    data[ 7622] = -'sd53187;
    data[ 7623] = -'sd44627;
    data[ 7624] =  'sd15293;
    data[ 7625] = -'sd56790;
    data[ 7626] = -'sd69848;
    data[ 7627] =  'sd2587;
    data[ 7628] =  'sd18109;
    data[ 7629] = -'sd37078;
    data[ 7630] =  'sd68136;
    data[ 7631] = -'sd14571;
    data[ 7632] =  'sd61844;
    data[ 7633] = -'sd58615;
    data[ 7634] =  'sd81218;
    data[ 7635] =  'sd77003;
    data[ 7636] =  'sd47498;
    data[ 7637] =  'sd4804;
    data[ 7638] =  'sd33628;
    data[ 7639] =  'sd71555;
    data[ 7640] =  'sd9362;
    data[ 7641] =  'sd65534;
    data[ 7642] = -'sd32785;
    data[ 7643] = -'sd65654;
    data[ 7644] =  'sd31945;
    data[ 7645] =  'sd59774;
    data[ 7646] = -'sd73105;
    data[ 7647] = -'sd20212;
    data[ 7648] =  'sd22357;
    data[ 7649] = -'sd7342;
    data[ 7650] = -'sd51394;
    data[ 7651] = -'sd32076;
    data[ 7652] = -'sd60691;
    data[ 7653] =  'sd66686;
    data[ 7654] = -'sd24721;
    data[ 7655] = -'sd9206;
    data[ 7656] = -'sd64442;
    data[ 7657] =  'sd40429;
    data[ 7658] = -'sd44679;
    data[ 7659] =  'sd14929;
    data[ 7660] = -'sd59338;
    data[ 7661] =  'sd76157;
    data[ 7662] =  'sd41576;
    data[ 7663] = -'sd36650;
    data[ 7664] =  'sd71132;
    data[ 7665] =  'sd6401;
    data[ 7666] =  'sd44807;
    data[ 7667] = -'sd14033;
    data[ 7668] =  'sd65610;
    data[ 7669] = -'sd32253;
    data[ 7670] = -'sd61930;
    data[ 7671] =  'sd58013;
    data[ 7672] =  'sd78409;
    data[ 7673] =  'sd57340;
    data[ 7674] =  'sd73698;
    data[ 7675] =  'sd24363;
    data[ 7676] =  'sd6700;
    data[ 7677] =  'sd46900;
    data[ 7678] =  'sd618;
    data[ 7679] =  'sd4326;
    data[ 7680] =  'sd30282;
    data[ 7681] =  'sd48133;
    data[ 7682] =  'sd9249;
    data[ 7683] =  'sd64743;
    data[ 7684] = -'sd38322;
    data[ 7685] =  'sd59428;
    data[ 7686] = -'sd75527;
    data[ 7687] = -'sd37166;
    data[ 7688] =  'sd67520;
    data[ 7689] = -'sd18883;
    data[ 7690] =  'sd31660;
    data[ 7691] =  'sd57779;
    data[ 7692] =  'sd76771;
    data[ 7693] =  'sd45874;
    data[ 7694] = -'sd6564;
    data[ 7695] = -'sd45948;
    data[ 7696] =  'sd6046;
    data[ 7697] =  'sd42322;
    data[ 7698] = -'sd31428;
    data[ 7699] = -'sd56155;
    data[ 7700] = -'sd65403;
    data[ 7701] =  'sd33702;
    data[ 7702] =  'sd72073;
    data[ 7703] =  'sd12988;
    data[ 7704] = -'sd72925;
    data[ 7705] = -'sd18952;
    data[ 7706] =  'sd31177;
    data[ 7707] =  'sd54398;
    data[ 7708] =  'sd53104;
    data[ 7709] =  'sd44046;
    data[ 7710] = -'sd19360;
    data[ 7711] =  'sd28321;
    data[ 7712] =  'sd34406;
    data[ 7713] =  'sd77001;
    data[ 7714] =  'sd47484;
    data[ 7715] =  'sd4706;
    data[ 7716] =  'sd32942;
    data[ 7717] =  'sd66753;
    data[ 7718] = -'sd24252;
    data[ 7719] = -'sd5923;
    data[ 7720] = -'sd41461;
    data[ 7721] =  'sd37455;
    data[ 7722] = -'sd65497;
    data[ 7723] =  'sd33044;
    data[ 7724] =  'sd67467;
    data[ 7725] = -'sd19254;
    data[ 7726] =  'sd29063;
    data[ 7727] =  'sd39600;
    data[ 7728] = -'sd50482;
    data[ 7729] = -'sd25692;
    data[ 7730] = -'sd16003;
    data[ 7731] =  'sd51820;
    data[ 7732] =  'sd35058;
    data[ 7733] =  'sd81565;
    data[ 7734] =  'sd79432;
    data[ 7735] =  'sd64501;
    data[ 7736] = -'sd40016;
    data[ 7737] =  'sd47570;
    data[ 7738] =  'sd5308;
    data[ 7739] =  'sd37156;
    data[ 7740] = -'sd67590;
    data[ 7741] =  'sd18393;
    data[ 7742] = -'sd35090;
    data[ 7743] = -'sd81789;
    data[ 7744] = -'sd81000;
    data[ 7745] = -'sd75477;
    data[ 7746] = -'sd36816;
    data[ 7747] =  'sd69970;
    data[ 7748] = -'sd1733;
    data[ 7749] = -'sd12131;
    data[ 7750] =  'sd78924;
    data[ 7751] =  'sd60945;
    data[ 7752] = -'sd64908;
    data[ 7753] =  'sd37167;
    data[ 7754] = -'sd67513;
    data[ 7755] =  'sd18932;
    data[ 7756] = -'sd31317;
    data[ 7757] = -'sd55378;
    data[ 7758] = -'sd59964;
    data[ 7759] =  'sd71775;
    data[ 7760] =  'sd10902;
    data[ 7761] =  'sd76314;
    data[ 7762] =  'sd42675;
    data[ 7763] = -'sd28957;
    data[ 7764] = -'sd38858;
    data[ 7765] =  'sd55676;
    data[ 7766] =  'sd62050;
    data[ 7767] = -'sd57173;
    data[ 7768] = -'sd72529;
    data[ 7769] = -'sd16180;
    data[ 7770] =  'sd50581;
    data[ 7771] =  'sd26385;
    data[ 7772] =  'sd20854;
    data[ 7773] = -'sd17863;
    data[ 7774] =  'sd38800;
    data[ 7775] = -'sd56082;
    data[ 7776] = -'sd64892;
    data[ 7777] =  'sd37279;
    data[ 7778] = -'sd66729;
    data[ 7779] =  'sd24420;
    data[ 7780] =  'sd7099;
    data[ 7781] =  'sd49693;
    data[ 7782] =  'sd20169;
    data[ 7783] = -'sd22658;
    data[ 7784] =  'sd5235;
    data[ 7785] =  'sd36645;
    data[ 7786] = -'sd71167;
    data[ 7787] = -'sd6646;
    data[ 7788] = -'sd46522;
    data[ 7789] =  'sd2028;
    data[ 7790] =  'sd14196;
    data[ 7791] = -'sd64469;
    data[ 7792] =  'sd40240;
    data[ 7793] = -'sd46002;
    data[ 7794] =  'sd5668;
    data[ 7795] =  'sd39676;
    data[ 7796] = -'sd49950;
    data[ 7797] = -'sd21968;
    data[ 7798] =  'sd10065;
    data[ 7799] =  'sd70455;
    data[ 7800] =  'sd1662;
    data[ 7801] =  'sd11634;
    data[ 7802] =  'sd81438;
    data[ 7803] =  'sd78543;
    data[ 7804] =  'sd58278;
    data[ 7805] =  'sd80264;
    data[ 7806] =  'sd70325;
    data[ 7807] =  'sd752;
    data[ 7808] =  'sd5264;
    data[ 7809] =  'sd36848;
    data[ 7810] = -'sd69746;
    data[ 7811] =  'sd3301;
    data[ 7812] =  'sd23107;
    data[ 7813] = -'sd2092;
    data[ 7814] = -'sd14644;
    data[ 7815] =  'sd61333;
    data[ 7816] = -'sd62192;
    data[ 7817] =  'sd56179;
    data[ 7818] =  'sd65571;
    data[ 7819] = -'sd32526;
    data[ 7820] = -'sd63841;
    data[ 7821] =  'sd44636;
    data[ 7822] = -'sd15230;
    data[ 7823] =  'sd57231;
    data[ 7824] =  'sd72935;
    data[ 7825] =  'sd19022;
    data[ 7826] = -'sd30687;
    data[ 7827] = -'sd50968;
    data[ 7828] = -'sd29094;
    data[ 7829] = -'sd39817;
    data[ 7830] =  'sd48963;
    data[ 7831] =  'sd15059;
    data[ 7832] = -'sd58428;
    data[ 7833] = -'sd81314;
    data[ 7834] = -'sd77675;
    data[ 7835] = -'sd52202;
    data[ 7836] = -'sd37732;
    data[ 7837] =  'sd63558;
    data[ 7838] = -'sd46617;
    data[ 7839] =  'sd1363;
    data[ 7840] =  'sd9541;
    data[ 7841] =  'sd66787;
    data[ 7842] = -'sd24014;
    data[ 7843] = -'sd4257;
    data[ 7844] = -'sd29799;
    data[ 7845] = -'sd44752;
    data[ 7846] =  'sd14418;
    data[ 7847] = -'sd62915;
    data[ 7848] =  'sd51118;
    data[ 7849] =  'sd30144;
    data[ 7850] =  'sd47167;
    data[ 7851] =  'sd2487;
    data[ 7852] =  'sd17409;
    data[ 7853] = -'sd41978;
    data[ 7854] =  'sd33836;
    data[ 7855] =  'sd73011;
    data[ 7856] =  'sd19554;
    data[ 7857] = -'sd26963;
    data[ 7858] = -'sd24900;
    data[ 7859] = -'sd10459;
    data[ 7860] = -'sd73213;
    data[ 7861] = -'sd20968;
    data[ 7862] =  'sd17065;
    data[ 7863] = -'sd44386;
    data[ 7864] =  'sd16980;
    data[ 7865] = -'sd44981;
    data[ 7866] =  'sd12815;
    data[ 7867] = -'sd74136;
    data[ 7868] = -'sd27429;
    data[ 7869] = -'sd28162;
    data[ 7870] = -'sd33293;
    data[ 7871] = -'sd69210;
    data[ 7872] =  'sd7053;
    data[ 7873] =  'sd49371;
    data[ 7874] =  'sd17915;
    data[ 7875] = -'sd38436;
    data[ 7876] =  'sd58630;
    data[ 7877] = -'sd81113;
    data[ 7878] = -'sd76268;
    data[ 7879] = -'sd42353;
    data[ 7880] =  'sd31211;
    data[ 7881] =  'sd54636;
    data[ 7882] =  'sd54770;
    data[ 7883] =  'sd55708;
    data[ 7884] =  'sd62274;
    data[ 7885] = -'sd55605;
    data[ 7886] = -'sd61553;
    data[ 7887] =  'sd60652;
    data[ 7888] = -'sd66959;
    data[ 7889] =  'sd22810;
    data[ 7890] = -'sd4171;
    data[ 7891] = -'sd29197;
    data[ 7892] = -'sd40538;
    data[ 7893] =  'sd43916;
    data[ 7894] = -'sd20270;
    data[ 7895] =  'sd21951;
    data[ 7896] = -'sd10184;
    data[ 7897] = -'sd71288;
    data[ 7898] = -'sd7493;
    data[ 7899] = -'sd52451;
    data[ 7900] = -'sd39475;
    data[ 7901] =  'sd51357;
    data[ 7902] =  'sd31817;
    data[ 7903] =  'sd58878;
    data[ 7904] = -'sd79377;
    data[ 7905] = -'sd64116;
    data[ 7906] =  'sd42711;
    data[ 7907] = -'sd28705;
    data[ 7908] = -'sd37094;
    data[ 7909] =  'sd68024;
    data[ 7910] = -'sd15355;
    data[ 7911] =  'sd56356;
    data[ 7912] =  'sd66810;
    data[ 7913] = -'sd23853;
    data[ 7914] = -'sd3130;
    data[ 7915] = -'sd21910;
    data[ 7916] =  'sd10471;
    data[ 7917] =  'sd73297;
    data[ 7918] =  'sd21556;
    data[ 7919] = -'sd12949;
    data[ 7920] =  'sd73198;
    data[ 7921] =  'sd20863;
    data[ 7922] = -'sd17800;
    data[ 7923] =  'sd39241;
    data[ 7924] = -'sd52995;
    data[ 7925] = -'sd43283;
    data[ 7926] =  'sd24701;
    data[ 7927] =  'sd9066;
    data[ 7928] =  'sd63462;
    data[ 7929] = -'sd47289;
    data[ 7930] = -'sd3341;
    data[ 7931] = -'sd23387;
    data[ 7932] =  'sd132;
    data[ 7933] =  'sd924;
    data[ 7934] =  'sd6468;
    data[ 7935] =  'sd45276;
    data[ 7936] = -'sd10750;
    data[ 7937] = -'sd75250;
    data[ 7938] = -'sd35227;
    data[ 7939] =  'sd81093;
    data[ 7940] =  'sd76128;
    data[ 7941] =  'sd41373;
    data[ 7942] = -'sd38071;
    data[ 7943] =  'sd61185;
    data[ 7944] = -'sd63228;
    data[ 7945] =  'sd48927;
    data[ 7946] =  'sd14807;
    data[ 7947] = -'sd60192;
    data[ 7948] =  'sd70179;
    data[ 7949] = -'sd270;
    data[ 7950] = -'sd1890;
    data[ 7951] = -'sd13230;
    data[ 7952] =  'sd71231;
    data[ 7953] =  'sd7094;
    data[ 7954] =  'sd49658;
    data[ 7955] =  'sd19924;
    data[ 7956] = -'sd24373;
    data[ 7957] = -'sd6770;
    data[ 7958] = -'sd47390;
    data[ 7959] = -'sd4048;
    data[ 7960] = -'sd28336;
    data[ 7961] = -'sd34511;
    data[ 7962] = -'sd77736;
    data[ 7963] = -'sd52629;
    data[ 7964] = -'sd40721;
    data[ 7965] =  'sd42635;
    data[ 7966] = -'sd29237;
    data[ 7967] = -'sd40818;
    data[ 7968] =  'sd41956;
    data[ 7969] = -'sd33990;
    data[ 7970] = -'sd74089;
    data[ 7971] = -'sd27100;
    data[ 7972] = -'sd25859;
    data[ 7973] = -'sd17172;
    data[ 7974] =  'sd43637;
    data[ 7975] = -'sd22223;
    data[ 7976] =  'sd8280;
    data[ 7977] =  'sd57960;
    data[ 7978] =  'sd78038;
    data[ 7979] =  'sd54743;
    data[ 7980] =  'sd55519;
    data[ 7981] =  'sd60951;
    data[ 7982] = -'sd64866;
    data[ 7983] =  'sd37461;
    data[ 7984] = -'sd65455;
    data[ 7985] =  'sd33338;
    data[ 7986] =  'sd69525;
    data[ 7987] = -'sd4848;
    data[ 7988] = -'sd33936;
    data[ 7989] = -'sd73711;
    data[ 7990] = -'sd24454;
    data[ 7991] = -'sd7337;
    data[ 7992] = -'sd51359;
    data[ 7993] = -'sd31831;
    data[ 7994] = -'sd58976;
    data[ 7995] =  'sd78691;
    data[ 7996] =  'sd59314;
    data[ 7997] = -'sd76325;
    data[ 7998] = -'sd42752;
    data[ 7999] =  'sd28418;
    data[ 8000] =  'sd35085;
    data[ 8001] =  'sd81754;
    data[ 8002] =  'sd80755;
    data[ 8003] =  'sd73762;
    data[ 8004] =  'sd24811;
    data[ 8005] =  'sd9836;
    data[ 8006] =  'sd68852;
    data[ 8007] = -'sd9559;
    data[ 8008] = -'sd66913;
    data[ 8009] =  'sd23132;
    data[ 8010] = -'sd1917;
    data[ 8011] = -'sd13419;
    data[ 8012] =  'sd69908;
    data[ 8013] = -'sd2167;
    data[ 8014] = -'sd15169;
    data[ 8015] =  'sd57658;
    data[ 8016] =  'sd75924;
    data[ 8017] =  'sd39945;
    data[ 8018] = -'sd48067;
    data[ 8019] = -'sd8787;
    data[ 8020] = -'sd61509;
    data[ 8021] =  'sd60960;
    data[ 8022] = -'sd64803;
    data[ 8023] =  'sd37902;
    data[ 8024] = -'sd62368;
    data[ 8025] =  'sd54947;
    data[ 8026] =  'sd56947;
    data[ 8027] =  'sd70947;
    data[ 8028] =  'sd5106;
    data[ 8029] =  'sd35742;
    data[ 8030] = -'sd77488;
    data[ 8031] = -'sd50893;
    data[ 8032] = -'sd28569;
    data[ 8033] = -'sd36142;
    data[ 8034] =  'sd74688;
    data[ 8035] =  'sd31293;
    data[ 8036] =  'sd55210;
    data[ 8037] =  'sd58788;
    data[ 8038] = -'sd80007;
    data[ 8039] = -'sd68526;
    data[ 8040] =  'sd11841;
    data[ 8041] = -'sd80954;
    data[ 8042] = -'sd75155;
    data[ 8043] = -'sd34562;
    data[ 8044] = -'sd78093;
    data[ 8045] = -'sd55128;
    data[ 8046] = -'sd58214;
    data[ 8047] = -'sd79816;
    data[ 8048] = -'sd67189;
    data[ 8049] =  'sd21200;
    data[ 8050] = -'sd15441;
    data[ 8051] =  'sd55754;
    data[ 8052] =  'sd62596;
    data[ 8053] = -'sd53351;
    data[ 8054] = -'sd45775;
    data[ 8055] =  'sd7257;
    data[ 8056] =  'sd50799;
    data[ 8057] =  'sd27911;
    data[ 8058] =  'sd31536;
    data[ 8059] =  'sd56911;
    data[ 8060] =  'sd70695;
    data[ 8061] =  'sd3342;
    data[ 8062] =  'sd23394;
    data[ 8063] = -'sd83;
    data[ 8064] = -'sd581;
    data[ 8065] = -'sd4067;
    data[ 8066] = -'sd28469;
    data[ 8067] = -'sd35442;
    data[ 8068] =  'sd79588;
    data[ 8069] =  'sd65593;
    data[ 8070] = -'sd32372;
    data[ 8071] = -'sd62763;
    data[ 8072] =  'sd52182;
    data[ 8073] =  'sd37592;
    data[ 8074] = -'sd64538;
    data[ 8075] =  'sd39757;
    data[ 8076] = -'sd49383;
    data[ 8077] = -'sd17999;
    data[ 8078] =  'sd37848;
    data[ 8079] = -'sd62746;
    data[ 8080] =  'sd52301;
    data[ 8081] =  'sd38425;
    data[ 8082] = -'sd58707;
    data[ 8083] =  'sd80574;
    data[ 8084] =  'sd72495;
    data[ 8085] =  'sd15942;
    data[ 8086] = -'sd52247;
    data[ 8087] = -'sd38047;
    data[ 8088] =  'sd61353;
    data[ 8089] = -'sd62052;
    data[ 8090] =  'sd57159;
    data[ 8091] =  'sd72431;
    data[ 8092] =  'sd15494;
    data[ 8093] = -'sd55383;
    data[ 8094] = -'sd59999;
    data[ 8095] =  'sd71530;
    data[ 8096] =  'sd9187;
    data[ 8097] =  'sd64309;
    data[ 8098] = -'sd41360;
    data[ 8099] =  'sd38162;
    data[ 8100] = -'sd60548;
    data[ 8101] =  'sd67687;
    data[ 8102] = -'sd17714;
    data[ 8103] =  'sd39843;
    data[ 8104] = -'sd48781;
    data[ 8105] = -'sd13785;
    data[ 8106] =  'sd67346;
    data[ 8107] = -'sd20101;
    data[ 8108] =  'sd23134;
    data[ 8109] = -'sd1903;
    data[ 8110] = -'sd13321;
    data[ 8111] =  'sd70594;
    data[ 8112] =  'sd2635;
    data[ 8113] =  'sd18445;
    data[ 8114] = -'sd34726;
    data[ 8115] = -'sd79241;
    data[ 8116] = -'sd63164;
    data[ 8117] =  'sd49375;
    data[ 8118] =  'sd17943;
    data[ 8119] = -'sd38240;
    data[ 8120] =  'sd60002;
    data[ 8121] = -'sd71509;
    data[ 8122] = -'sd9040;
    data[ 8123] = -'sd63280;
    data[ 8124] =  'sd48563;
    data[ 8125] =  'sd12259;
    data[ 8126] = -'sd78028;
    data[ 8127] = -'sd54673;
    data[ 8128] = -'sd55029;
    data[ 8129] = -'sd57521;
    data[ 8130] = -'sd74965;
    data[ 8131] = -'sd33232;
    data[ 8132] = -'sd68783;
    data[ 8133] =  'sd10042;
    data[ 8134] =  'sd70294;
    data[ 8135] =  'sd535;
    data[ 8136] =  'sd3745;
    data[ 8137] =  'sd26215;
    data[ 8138] =  'sd19664;
    data[ 8139] = -'sd26193;
    data[ 8140] = -'sd19510;
    data[ 8141] =  'sd27271;
    data[ 8142] =  'sd27056;
    data[ 8143] =  'sd25551;
    data[ 8144] =  'sd15016;
    data[ 8145] = -'sd58729;
    data[ 8146] =  'sd80420;
    data[ 8147] =  'sd71417;
    data[ 8148] =  'sd8396;
    data[ 8149] =  'sd58772;
    data[ 8150] = -'sd80119;
    data[ 8151] = -'sd69310;
    data[ 8152] =  'sd6353;
    data[ 8153] =  'sd44471;
    data[ 8154] = -'sd16385;
    data[ 8155] =  'sd49146;
    data[ 8156] =  'sd16340;
    data[ 8157] = -'sd49461;
    data[ 8158] = -'sd18545;
    data[ 8159] =  'sd34026;
    data[ 8160] =  'sd74341;
    data[ 8161] =  'sd28864;
    data[ 8162] =  'sd38207;
    data[ 8163] = -'sd60233;
    data[ 8164] =  'sd69892;
    data[ 8165] = -'sd2279;
    data[ 8166] = -'sd15953;
    data[ 8167] =  'sd52170;
    data[ 8168] =  'sd37508;
    data[ 8169] = -'sd65126;
    data[ 8170] =  'sd35641;
    data[ 8171] = -'sd78195;
    data[ 8172] = -'sd55842;
    data[ 8173] = -'sd63212;
    data[ 8174] =  'sd49039;
    data[ 8175] =  'sd15591;
    data[ 8176] = -'sd54704;
    data[ 8177] = -'sd55246;
    data[ 8178] = -'sd59040;
    data[ 8179] =  'sd78243;
    data[ 8180] =  'sd56178;
    data[ 8181] =  'sd65564;
    data[ 8182] = -'sd32575;
    data[ 8183] = -'sd64184;
    data[ 8184] =  'sd42235;
    data[ 8185] = -'sd32037;
    data[ 8186] = -'sd60418;
    data[ 8187] =  'sd68597;
    data[ 8188] = -'sd11344;
    data[ 8189] = -'sd79408;
    data[ 8190] = -'sd64333;
    data[ 8191] =  'sd41192;
    data[ 8192] = -'sd39338;
    data[ 8193] =  'sd52316;
    data[ 8194] =  'sd38530;
    data[ 8195] = -'sd57972;
    data[ 8196] = -'sd78122;
    data[ 8197] = -'sd55331;
    data[ 8198] = -'sd59635;
    data[ 8199] =  'sd74078;
    data[ 8200] =  'sd27023;
    data[ 8201] =  'sd25320;
    data[ 8202] =  'sd13399;
    data[ 8203] = -'sd70048;
    data[ 8204] =  'sd1187;
    data[ 8205] =  'sd8309;
    data[ 8206] =  'sd58163;
    data[ 8207] =  'sd79459;
    data[ 8208] =  'sd64690;
    data[ 8209] = -'sd38693;
    data[ 8210] =  'sd56831;
    data[ 8211] =  'sd70135;
    data[ 8212] = -'sd578;
    data[ 8213] = -'sd4046;
    data[ 8214] = -'sd28322;
    data[ 8215] = -'sd34413;
    data[ 8216] = -'sd77050;
    data[ 8217] = -'sd47827;
    data[ 8218] = -'sd7107;
    data[ 8219] = -'sd49749;
    data[ 8220] = -'sd20561;
    data[ 8221] =  'sd19914;
    data[ 8222] = -'sd24443;
    data[ 8223] = -'sd7260;
    data[ 8224] = -'sd50820;
    data[ 8225] = -'sd28058;
    data[ 8226] = -'sd32565;
    data[ 8227] = -'sd64114;
    data[ 8228] =  'sd42725;
    data[ 8229] = -'sd28607;
    data[ 8230] = -'sd36408;
    data[ 8231] =  'sd72826;
    data[ 8232] =  'sd18259;
    data[ 8233] = -'sd36028;
    data[ 8234] =  'sd75486;
    data[ 8235] =  'sd36879;
    data[ 8236] = -'sd69529;
    data[ 8237] =  'sd4820;
    data[ 8238] =  'sd33740;
    data[ 8239] =  'sd72339;
    data[ 8240] =  'sd14850;
    data[ 8241] = -'sd59891;
    data[ 8242] =  'sd72286;
    data[ 8243] =  'sd14479;
    data[ 8244] = -'sd62488;
    data[ 8245] =  'sd54107;
    data[ 8246] =  'sd51067;
    data[ 8247] =  'sd29787;
    data[ 8248] =  'sd44668;
    data[ 8249] = -'sd15006;
    data[ 8250] =  'sd58799;
    data[ 8251] = -'sd79930;
    data[ 8252] = -'sd67987;
    data[ 8253] =  'sd15614;
    data[ 8254] = -'sd54543;
    data[ 8255] = -'sd54119;
    data[ 8256] = -'sd51151;
    data[ 8257] = -'sd30375;
    data[ 8258] = -'sd48784;
    data[ 8259] = -'sd13806;
    data[ 8260] =  'sd67199;
    data[ 8261] = -'sd21130;
    data[ 8262] =  'sd15931;
    data[ 8263] = -'sd52324;
    data[ 8264] = -'sd38586;
    data[ 8265] =  'sd57580;
    data[ 8266] =  'sd75378;
    data[ 8267] =  'sd36123;
    data[ 8268] = -'sd74821;
    data[ 8269] = -'sd32224;
    data[ 8270] = -'sd61727;
    data[ 8271] =  'sd59434;
    data[ 8272] = -'sd75485;
    data[ 8273] = -'sd36872;
    data[ 8274] =  'sd69578;
    data[ 8275] = -'sd4477;
    data[ 8276] = -'sd31339;
    data[ 8277] = -'sd55532;
    data[ 8278] = -'sd61042;
    data[ 8279] =  'sd64229;
    data[ 8280] = -'sd41920;
    data[ 8281] =  'sd34242;
    data[ 8282] =  'sd75853;
    data[ 8283] =  'sd39448;
    data[ 8284] = -'sd51546;
    data[ 8285] = -'sd33140;
    data[ 8286] = -'sd68139;
    data[ 8287] =  'sd14550;
    data[ 8288] = -'sd61991;
    data[ 8289] =  'sd57586;
    data[ 8290] =  'sd75420;
    data[ 8291] =  'sd36417;
    data[ 8292] = -'sd72763;
    data[ 8293] = -'sd17818;
    data[ 8294] =  'sd39115;
    data[ 8295] = -'sd53877;
    data[ 8296] = -'sd49457;
    data[ 8297] = -'sd18517;
    data[ 8298] =  'sd34222;
    data[ 8299] =  'sd75713;
    data[ 8300] =  'sd38468;
    data[ 8301] = -'sd58406;
    data[ 8302] = -'sd81160;
    data[ 8303] = -'sd76597;
    data[ 8304] = -'sd44656;
    data[ 8305] =  'sd15090;
    data[ 8306] = -'sd58211;
    data[ 8307] = -'sd79795;
    data[ 8308] = -'sd67042;
    data[ 8309] =  'sd22229;
    data[ 8310] = -'sd8238;
    data[ 8311] = -'sd57666;
    data[ 8312] = -'sd75980;
    data[ 8313] = -'sd40337;
    data[ 8314] =  'sd45323;
    data[ 8315] = -'sd10421;
    data[ 8316] = -'sd72947;
    data[ 8317] = -'sd19106;
    data[ 8318] =  'sd30099;
    data[ 8319] =  'sd46852;
    data[ 8320] =  'sd282;
    data[ 8321] =  'sd1974;
    data[ 8322] =  'sd13818;
    data[ 8323] = -'sd67115;
    data[ 8324] =  'sd21718;
    data[ 8325] = -'sd11815;
    data[ 8326] =  'sd81136;
    data[ 8327] =  'sd76429;
    data[ 8328] =  'sd43480;
    data[ 8329] = -'sd23322;
    data[ 8330] =  'sd587;
    data[ 8331] =  'sd4109;
    data[ 8332] =  'sd28763;
    data[ 8333] =  'sd37500;
    data[ 8334] = -'sd65182;
    data[ 8335] =  'sd35249;
    data[ 8336] = -'sd80939;
    data[ 8337] = -'sd75050;
    data[ 8338] = -'sd33827;
    data[ 8339] = -'sd72948;
    data[ 8340] = -'sd19113;
    data[ 8341] =  'sd30050;
    data[ 8342] =  'sd46509;
    data[ 8343] = -'sd2119;
    data[ 8344] = -'sd14833;
    data[ 8345] =  'sd60010;
    data[ 8346] = -'sd71453;
    data[ 8347] = -'sd8648;
    data[ 8348] = -'sd60536;
    data[ 8349] =  'sd67771;
    data[ 8350] = -'sd17126;
    data[ 8351] =  'sd43959;
    data[ 8352] = -'sd19969;
    data[ 8353] =  'sd24058;
    data[ 8354] =  'sd4565;
    data[ 8355] =  'sd31955;
    data[ 8356] =  'sd59844;
    data[ 8357] = -'sd72615;
    data[ 8358] = -'sd16782;
    data[ 8359] =  'sd46367;
    data[ 8360] = -'sd3113;
    data[ 8361] = -'sd21791;
    data[ 8362] =  'sd11304;
    data[ 8363] =  'sd79128;
    data[ 8364] =  'sd62373;
    data[ 8365] = -'sd54912;
    data[ 8366] = -'sd56702;
    data[ 8367] = -'sd69232;
    data[ 8368] =  'sd6899;
    data[ 8369] =  'sd48293;
    data[ 8370] =  'sd10369;
    data[ 8371] =  'sd72583;
    data[ 8372] =  'sd16558;
    data[ 8373] = -'sd47935;
    data[ 8374] = -'sd7863;
    data[ 8375] = -'sd55041;
    data[ 8376] = -'sd57605;
    data[ 8377] = -'sd75553;
    data[ 8378] = -'sd37348;
    data[ 8379] =  'sd66246;
    data[ 8380] = -'sd27801;
    data[ 8381] = -'sd30766;
    data[ 8382] = -'sd51521;
    data[ 8383] = -'sd32965;
    data[ 8384] = -'sd66914;
    data[ 8385] =  'sd23125;
    data[ 8386] = -'sd1966;
    data[ 8387] = -'sd13762;
    data[ 8388] =  'sd67507;
    data[ 8389] = -'sd18974;
    data[ 8390] =  'sd31023;
    data[ 8391] =  'sd53320;
    data[ 8392] =  'sd45558;
    data[ 8393] = -'sd8776;
    data[ 8394] = -'sd61432;
    data[ 8395] =  'sd61499;
    data[ 8396] = -'sd61030;
    data[ 8397] =  'sd64313;
    data[ 8398] = -'sd41332;
    data[ 8399] =  'sd38358;
    data[ 8400] = -'sd59176;
    data[ 8401] =  'sd77291;
    data[ 8402] =  'sd49514;
    data[ 8403] =  'sd18916;
    data[ 8404] = -'sd31429;
    data[ 8405] = -'sd56162;
    data[ 8406] = -'sd65452;
    data[ 8407] =  'sd33359;
    data[ 8408] =  'sd69672;
    data[ 8409] = -'sd3819;
    data[ 8410] = -'sd26733;
    data[ 8411] = -'sd23290;
    data[ 8412] =  'sd811;
    data[ 8413] =  'sd5677;
    data[ 8414] =  'sd39739;
    data[ 8415] = -'sd49509;
    data[ 8416] = -'sd18881;
    data[ 8417] =  'sd31674;
    data[ 8418] =  'sd57877;
    data[ 8419] =  'sd77457;
    data[ 8420] =  'sd50676;
    data[ 8421] =  'sd27050;
    data[ 8422] =  'sd25509;
    data[ 8423] =  'sd14722;
    data[ 8424] = -'sd60787;
    data[ 8425] =  'sd66014;
    data[ 8426] = -'sd29425;
    data[ 8427] = -'sd42134;
    data[ 8428] =  'sd32744;
    data[ 8429] =  'sd65367;
    data[ 8430] = -'sd33954;
    data[ 8431] = -'sd73837;
    data[ 8432] = -'sd25336;
    data[ 8433] = -'sd13511;
    data[ 8434] =  'sd69264;
    data[ 8435] = -'sd6675;
    data[ 8436] = -'sd46725;
    data[ 8437] =  'sd607;
    data[ 8438] =  'sd4249;
    data[ 8439] =  'sd29743;
    data[ 8440] =  'sd44360;
    data[ 8441] = -'sd17162;
    data[ 8442] =  'sd43707;
    data[ 8443] = -'sd21733;
    data[ 8444] =  'sd11710;
    data[ 8445] = -'sd81871;
    data[ 8446] = -'sd81574;
    data[ 8447] = -'sd79495;
    data[ 8448] = -'sd64942;
    data[ 8449] =  'sd36929;
    data[ 8450] = -'sd69179;
    data[ 8451] =  'sd7270;
    data[ 8452] =  'sd50890;
    data[ 8453] =  'sd28548;
    data[ 8454] =  'sd35995;
    data[ 8455] = -'sd75717;
    data[ 8456] = -'sd38496;
    data[ 8457] =  'sd58210;
    data[ 8458] =  'sd79788;
    data[ 8459] =  'sd66993;
    data[ 8460] = -'sd22572;
    data[ 8461] =  'sd5837;
    data[ 8462] =  'sd40859;
    data[ 8463] = -'sd41669;
    data[ 8464] =  'sd35999;
    data[ 8465] = -'sd75689;
    data[ 8466] = -'sd38300;
    data[ 8467] =  'sd59582;
    data[ 8468] = -'sd74449;
    data[ 8469] = -'sd29620;
    data[ 8470] = -'sd43499;
    data[ 8471] =  'sd23189;
    data[ 8472] = -'sd1518;
    data[ 8473] = -'sd10626;
    data[ 8474] = -'sd74382;
    data[ 8475] = -'sd29151;
    data[ 8476] = -'sd40216;
    data[ 8477] =  'sd46170;
    data[ 8478] = -'sd4492;
    data[ 8479] = -'sd31444;
    data[ 8480] = -'sd56267;
    data[ 8481] = -'sd66187;
    data[ 8482] =  'sd28214;
    data[ 8483] =  'sd33657;
    data[ 8484] =  'sd71758;
    data[ 8485] =  'sd10783;
    data[ 8486] =  'sd75481;
    data[ 8487] =  'sd36844;
    data[ 8488] = -'sd69774;
    data[ 8489] =  'sd3105;
    data[ 8490] =  'sd21735;
    data[ 8491] = -'sd11696;
    data[ 8492] = -'sd81872;
    data[ 8493] = -'sd81581;
    data[ 8494] = -'sd79544;
    data[ 8495] = -'sd65285;
    data[ 8496] =  'sd34528;
    data[ 8497] =  'sd77855;
    data[ 8498] =  'sd53462;
    data[ 8499] =  'sd46552;
    data[ 8500] = -'sd1818;
    data[ 8501] = -'sd12726;
    data[ 8502] =  'sd74759;
    data[ 8503] =  'sd31790;
    data[ 8504] =  'sd58689;
    data[ 8505] = -'sd80700;
    data[ 8506] = -'sd73377;
    data[ 8507] = -'sd22116;
    data[ 8508] =  'sd9029;
    data[ 8509] =  'sd63203;
    data[ 8510] = -'sd49102;
    data[ 8511] = -'sd16032;
    data[ 8512] =  'sd51617;
    data[ 8513] =  'sd33637;
    data[ 8514] =  'sd71618;
    data[ 8515] =  'sd9803;
    data[ 8516] =  'sd68621;
    data[ 8517] = -'sd11176;
    data[ 8518] = -'sd78232;
    data[ 8519] = -'sd56101;
    data[ 8520] = -'sd65025;
    data[ 8521] =  'sd36348;
    data[ 8522] = -'sd73246;
    data[ 8523] = -'sd21199;
    data[ 8524] =  'sd15448;
    data[ 8525] = -'sd55705;
    data[ 8526] = -'sd62253;
    data[ 8527] =  'sd55752;
    data[ 8528] =  'sd62582;
    data[ 8529] = -'sd53449;
    data[ 8530] = -'sd46461;
    data[ 8531] =  'sd2455;
    data[ 8532] =  'sd17185;
    data[ 8533] = -'sd43546;
    data[ 8534] =  'sd22860;
    data[ 8535] = -'sd3821;
    data[ 8536] = -'sd26747;
    data[ 8537] = -'sd23388;
    data[ 8538] =  'sd125;
    data[ 8539] =  'sd875;
    data[ 8540] =  'sd6125;
    data[ 8541] =  'sd42875;
    data[ 8542] = -'sd27557;
    data[ 8543] = -'sd29058;
    data[ 8544] = -'sd39565;
    data[ 8545] =  'sd50727;
    data[ 8546] =  'sd27407;
    data[ 8547] =  'sd28008;
    data[ 8548] =  'sd32215;
    data[ 8549] =  'sd61664;
    data[ 8550] = -'sd59875;
    data[ 8551] =  'sd72398;
    data[ 8552] =  'sd15263;
    data[ 8553] = -'sd57000;
    data[ 8554] = -'sd71318;
    data[ 8555] = -'sd7703;
    data[ 8556] = -'sd53921;
    data[ 8557] = -'sd49765;
    data[ 8558] = -'sd20673;
    data[ 8559] =  'sd19130;
    data[ 8560] = -'sd29931;
    data[ 8561] = -'sd45676;
    data[ 8562] =  'sd7950;
    data[ 8563] =  'sd55650;
    data[ 8564] =  'sd61868;
    data[ 8565] = -'sd58447;
    data[ 8566] = -'sd81447;
    data[ 8567] = -'sd78606;
    data[ 8568] = -'sd58719;
    data[ 8569] =  'sd80490;
    data[ 8570] =  'sd71907;
    data[ 8571] =  'sd11826;
    data[ 8572] = -'sd81059;
    data[ 8573] = -'sd75890;
    data[ 8574] = -'sd39707;
    data[ 8575] =  'sd49733;
    data[ 8576] =  'sd20449;
    data[ 8577] = -'sd20698;
    data[ 8578] =  'sd18955;
    data[ 8579] = -'sd31156;
    data[ 8580] = -'sd54251;
    data[ 8581] = -'sd52075;
    data[ 8582] = -'sd36843;
    data[ 8583] =  'sd69781;
    data[ 8584] = -'sd3056;
    data[ 8585] = -'sd21392;
    data[ 8586] =  'sd14097;
    data[ 8587] = -'sd65162;
    data[ 8588] =  'sd35389;
    data[ 8589] = -'sd79959;
    data[ 8590] = -'sd68190;
    data[ 8591] =  'sd14193;
    data[ 8592] = -'sd64490;
    data[ 8593] =  'sd40093;
    data[ 8594] = -'sd47031;
    data[ 8595] = -'sd1535;
    data[ 8596] = -'sd10745;
    data[ 8597] = -'sd75215;
    data[ 8598] = -'sd34982;
    data[ 8599] = -'sd81033;
    data[ 8600] = -'sd75708;
    data[ 8601] = -'sd38433;
    data[ 8602] =  'sd58651;
    data[ 8603] = -'sd80966;
    data[ 8604] = -'sd75239;
    data[ 8605] = -'sd35150;
    data[ 8606] =  'sd81632;
    data[ 8607] =  'sd79901;
    data[ 8608] =  'sd67784;
    data[ 8609] = -'sd17035;
    data[ 8610] =  'sd44596;
    data[ 8611] = -'sd15510;
    data[ 8612] =  'sd55271;
    data[ 8613] =  'sd59215;
    data[ 8614] = -'sd77018;
    data[ 8615] = -'sd47603;
    data[ 8616] = -'sd5539;
    data[ 8617] = -'sd38773;
    data[ 8618] =  'sd56271;
    data[ 8619] =  'sd66215;
    data[ 8620] = -'sd28018;
    data[ 8621] = -'sd32285;
    data[ 8622] = -'sd62154;
    data[ 8623] =  'sd56445;
    data[ 8624] =  'sd67433;
    data[ 8625] = -'sd19492;
    data[ 8626] =  'sd27397;
    data[ 8627] =  'sd27938;
    data[ 8628] =  'sd31725;
    data[ 8629] =  'sd58234;
    data[ 8630] =  'sd79956;
    data[ 8631] =  'sd68169;
    data[ 8632] = -'sd14340;
    data[ 8633] =  'sd63461;
    data[ 8634] = -'sd47296;
    data[ 8635] = -'sd3390;
    data[ 8636] = -'sd23730;
    data[ 8637] = -'sd2269;
    data[ 8638] = -'sd15883;
    data[ 8639] =  'sd52660;
    data[ 8640] =  'sd40938;
    data[ 8641] = -'sd41116;
    data[ 8642] =  'sd39870;
    data[ 8643] = -'sd48592;
    data[ 8644] = -'sd12462;
    data[ 8645] =  'sd76607;
    data[ 8646] =  'sd44726;
    data[ 8647] = -'sd14600;
    data[ 8648] =  'sd61641;
    data[ 8649] = -'sd60036;
    data[ 8650] =  'sd71271;
    data[ 8651] =  'sd7374;
    data[ 8652] =  'sd51618;
    data[ 8653] =  'sd33644;
    data[ 8654] =  'sd71667;
    data[ 8655] =  'sd10146;
    data[ 8656] =  'sd71022;
    data[ 8657] =  'sd5631;
    data[ 8658] =  'sd39417;
    data[ 8659] = -'sd51763;
    data[ 8660] = -'sd34659;
    data[ 8661] = -'sd78772;
    data[ 8662] = -'sd59881;
    data[ 8663] =  'sd72356;
    data[ 8664] =  'sd14969;
    data[ 8665] = -'sd59058;
    data[ 8666] =  'sd78117;
    data[ 8667] =  'sd55296;
    data[ 8668] =  'sd59390;
    data[ 8669] = -'sd75793;
    data[ 8670] = -'sd39028;
    data[ 8671] =  'sd54486;
    data[ 8672] =  'sd53720;
    data[ 8673] =  'sd48358;
    data[ 8674] =  'sd10824;
    data[ 8675] =  'sd75768;
    data[ 8676] =  'sd38853;
    data[ 8677] = -'sd55711;
    data[ 8678] = -'sd62295;
    data[ 8679] =  'sd55458;
    data[ 8680] =  'sd60524;
    data[ 8681] = -'sd67855;
    data[ 8682] =  'sd16538;
    data[ 8683] = -'sd48075;
    data[ 8684] = -'sd8843;
    data[ 8685] = -'sd61901;
    data[ 8686] =  'sd58216;
    data[ 8687] =  'sd79830;
    data[ 8688] =  'sd67287;
    data[ 8689] = -'sd20514;
    data[ 8690] =  'sd20243;
    data[ 8691] = -'sd22140;
    data[ 8692] =  'sd8861;
    data[ 8693] =  'sd62027;
    data[ 8694] = -'sd57334;
    data[ 8695] = -'sd73656;
    data[ 8696] = -'sd24069;
    data[ 8697] = -'sd4642;
    data[ 8698] = -'sd32494;
    data[ 8699] = -'sd63617;
    data[ 8700] =  'sd46204;
    data[ 8701] = -'sd4254;
    data[ 8702] = -'sd29778;
    data[ 8703] = -'sd44605;
    data[ 8704] =  'sd15447;
    data[ 8705] = -'sd55712;
    data[ 8706] = -'sd62302;
    data[ 8707] =  'sd55409;
    data[ 8708] =  'sd60181;
    data[ 8709] = -'sd70256;
    data[ 8710] = -'sd269;
    data[ 8711] = -'sd1883;
    data[ 8712] = -'sd13181;
    data[ 8713] =  'sd71574;
    data[ 8714] =  'sd9495;
    data[ 8715] =  'sd66465;
    data[ 8716] = -'sd26268;
    data[ 8717] = -'sd20035;
    data[ 8718] =  'sd23596;
    data[ 8719] =  'sd1331;
    data[ 8720] =  'sd9317;
    data[ 8721] =  'sd65219;
    data[ 8722] = -'sd34990;
    data[ 8723] = -'sd81089;
    data[ 8724] = -'sd76100;
    data[ 8725] = -'sd41177;
    data[ 8726] =  'sd39443;
    data[ 8727] = -'sd51581;
    data[ 8728] = -'sd33385;
    data[ 8729] = -'sd69854;
    data[ 8730] =  'sd2545;
    data[ 8731] =  'sd17815;
    data[ 8732] = -'sd39136;
    data[ 8733] =  'sd53730;
    data[ 8734] =  'sd48428;
    data[ 8735] =  'sd11314;
    data[ 8736] =  'sd79198;
    data[ 8737] =  'sd62863;
    data[ 8738] = -'sd51482;
    data[ 8739] = -'sd32692;
    data[ 8740] = -'sd65003;
    data[ 8741] =  'sd36502;
    data[ 8742] = -'sd72168;
    data[ 8743] = -'sd13653;
    data[ 8744] =  'sd68270;
    data[ 8745] = -'sd13633;
    data[ 8746] =  'sd68410;
    data[ 8747] = -'sd12653;
    data[ 8748] =  'sd75270;
    data[ 8749] =  'sd35367;
    data[ 8750] = -'sd80113;
    data[ 8751] = -'sd69268;
    data[ 8752] =  'sd6647;
    data[ 8753] =  'sd46529;
    data[ 8754] = -'sd1979;
    data[ 8755] = -'sd13853;
    data[ 8756] =  'sd66870;
    data[ 8757] = -'sd23433;
    data[ 8758] = -'sd190;
    data[ 8759] = -'sd1330;
    data[ 8760] = -'sd9310;
    data[ 8761] = -'sd65170;
    data[ 8762] =  'sd35333;
    data[ 8763] = -'sd80351;
    data[ 8764] = -'sd70934;
    data[ 8765] = -'sd5015;
    data[ 8766] = -'sd35105;
    data[ 8767] = -'sd81894;
    data[ 8768] = -'sd81735;
    data[ 8769] = -'sd80622;
    data[ 8770] = -'sd72831;
    data[ 8771] = -'sd18294;
    data[ 8772] =  'sd35783;
    data[ 8773] = -'sd77201;
    data[ 8774] = -'sd48884;
    data[ 8775] = -'sd14506;
    data[ 8776] =  'sd62299;
    data[ 8777] = -'sd55430;
    data[ 8778] = -'sd60328;
    data[ 8779] =  'sd69227;
    data[ 8780] = -'sd6934;
    data[ 8781] = -'sd48538;
    data[ 8782] = -'sd12084;
    data[ 8783] =  'sd79253;
    data[ 8784] =  'sd63248;
    data[ 8785] = -'sd48787;
    data[ 8786] = -'sd13827;
    data[ 8787] =  'sd67052;
    data[ 8788] = -'sd22159;
    data[ 8789] =  'sd8728;
    data[ 8790] =  'sd61096;
    data[ 8791] = -'sd63851;
    data[ 8792] =  'sd44566;
    data[ 8793] = -'sd15720;
    data[ 8794] =  'sd53801;
    data[ 8795] =  'sd48925;
    data[ 8796] =  'sd14793;
    data[ 8797] = -'sd60290;
    data[ 8798] =  'sd69493;
    data[ 8799] = -'sd5072;
    data[ 8800] = -'sd35504;
    data[ 8801] =  'sd79154;
    data[ 8802] =  'sd62555;
    data[ 8803] = -'sd53638;
    data[ 8804] = -'sd47784;
    data[ 8805] = -'sd6806;
    data[ 8806] = -'sd47642;
    data[ 8807] = -'sd5812;
    data[ 8808] = -'sd40684;
    data[ 8809] =  'sd42894;
    data[ 8810] = -'sd27424;
    data[ 8811] = -'sd28127;
    data[ 8812] = -'sd33048;
    data[ 8813] = -'sd67495;
    data[ 8814] =  'sd19058;
    data[ 8815] = -'sd30435;
    data[ 8816] = -'sd49204;
    data[ 8817] = -'sd16746;
    data[ 8818] =  'sd46619;
    data[ 8819] = -'sd1349;
    data[ 8820] = -'sd9443;
    data[ 8821] = -'sd66101;
    data[ 8822] =  'sd28816;
    data[ 8823] =  'sd37871;
    data[ 8824] = -'sd62585;
    data[ 8825] =  'sd53428;
    data[ 8826] =  'sd46314;
    data[ 8827] = -'sd3484;
    data[ 8828] = -'sd24388;
    data[ 8829] = -'sd6875;
    data[ 8830] = -'sd48125;
    data[ 8831] = -'sd9193;
    data[ 8832] = -'sd64351;
    data[ 8833] =  'sd41066;
    data[ 8834] = -'sd40220;
    data[ 8835] =  'sd46142;
    data[ 8836] = -'sd4688;
    data[ 8837] = -'sd32816;
    data[ 8838] = -'sd65871;
    data[ 8839] =  'sd30426;
    data[ 8840] =  'sd49141;
    data[ 8841] =  'sd16305;
    data[ 8842] = -'sd49706;
    data[ 8843] = -'sd20260;
    data[ 8844] =  'sd22021;
    data[ 8845] = -'sd9694;
    data[ 8846] = -'sd67858;
    data[ 8847] =  'sd16517;
    data[ 8848] = -'sd48222;
    data[ 8849] = -'sd9872;
    data[ 8850] = -'sd69104;
    data[ 8851] =  'sd7795;
    data[ 8852] =  'sd54565;
    data[ 8853] =  'sd54273;
    data[ 8854] =  'sd52229;
    data[ 8855] =  'sd37921;
    data[ 8856] = -'sd62235;
    data[ 8857] =  'sd55878;
    data[ 8858] =  'sd63464;
    data[ 8859] = -'sd47275;
    data[ 8860] = -'sd3243;
    data[ 8861] = -'sd22701;
    data[ 8862] =  'sd4934;
    data[ 8863] =  'sd34538;
    data[ 8864] =  'sd77925;
    data[ 8865] =  'sd53952;
    data[ 8866] =  'sd49982;
    data[ 8867] =  'sd22192;
    data[ 8868] = -'sd8497;
    data[ 8869] = -'sd59479;
    data[ 8870] =  'sd75170;
    data[ 8871] =  'sd34667;
    data[ 8872] =  'sd78828;
    data[ 8873] =  'sd60273;
    data[ 8874] = -'sd69612;
    data[ 8875] =  'sd4239;
    data[ 8876] =  'sd29673;
    data[ 8877] =  'sd43870;
    data[ 8878] = -'sd20592;
    data[ 8879] =  'sd19697;
    data[ 8880] = -'sd25962;
    data[ 8881] = -'sd17893;
    data[ 8882] =  'sd38590;
    data[ 8883] = -'sd57552;
    data[ 8884] = -'sd75182;
    data[ 8885] = -'sd34751;
    data[ 8886] = -'sd79416;
    data[ 8887] = -'sd64389;
    data[ 8888] =  'sd40800;
    data[ 8889] = -'sd42082;
    data[ 8890] =  'sd33108;
    data[ 8891] =  'sd67915;
    data[ 8892] = -'sd16118;
    data[ 8893] =  'sd51015;
    data[ 8894] =  'sd29423;
    data[ 8895] =  'sd42120;
    data[ 8896] = -'sd32842;
    data[ 8897] = -'sd66053;
    data[ 8898] =  'sd29152;
    data[ 8899] =  'sd40223;
    data[ 8900] = -'sd46121;
    data[ 8901] =  'sd4835;
    data[ 8902] =  'sd33845;
    data[ 8903] =  'sd73074;
    data[ 8904] =  'sd19995;
    data[ 8905] = -'sd23876;
    data[ 8906] = -'sd3291;
    data[ 8907] = -'sd23037;
    data[ 8908] =  'sd2582;
    data[ 8909] =  'sd18074;
    data[ 8910] = -'sd37323;
    data[ 8911] =  'sd66421;
    data[ 8912] = -'sd26576;
    data[ 8913] = -'sd22191;
    data[ 8914] =  'sd8504;
    data[ 8915] =  'sd59528;
    data[ 8916] = -'sd74827;
    data[ 8917] = -'sd32266;
    data[ 8918] = -'sd62021;
    data[ 8919] =  'sd57376;
    data[ 8920] =  'sd73950;
    data[ 8921] =  'sd26127;
    data[ 8922] =  'sd19048;
    data[ 8923] = -'sd30505;
    data[ 8924] = -'sd49694;
    data[ 8925] = -'sd20176;
    data[ 8926] =  'sd22609;
    data[ 8927] = -'sd5578;
    data[ 8928] = -'sd39046;
    data[ 8929] =  'sd54360;
    data[ 8930] =  'sd52838;
    data[ 8931] =  'sd42184;
    data[ 8932] = -'sd32394;
    data[ 8933] = -'sd62917;
    data[ 8934] =  'sd51104;
    data[ 8935] =  'sd30046;
    data[ 8936] =  'sd46481;
    data[ 8937] = -'sd2315;
    data[ 8938] = -'sd16205;
    data[ 8939] =  'sd50406;
    data[ 8940] =  'sd25160;
    data[ 8941] =  'sd12279;
    data[ 8942] = -'sd77888;
    data[ 8943] = -'sd53693;
    data[ 8944] = -'sd48169;
    data[ 8945] = -'sd9501;
    data[ 8946] = -'sd66507;
    data[ 8947] =  'sd25974;
    data[ 8948] =  'sd17977;
    data[ 8949] = -'sd38002;
    data[ 8950] =  'sd61668;
    data[ 8951] = -'sd59847;
    data[ 8952] =  'sd72594;
    data[ 8953] =  'sd16635;
    data[ 8954] = -'sd47396;
    data[ 8955] = -'sd4090;
    data[ 8956] = -'sd28630;
    data[ 8957] = -'sd36569;
    data[ 8958] =  'sd71699;
    data[ 8959] =  'sd10370;
    data[ 8960] =  'sd72590;
    data[ 8961] =  'sd16607;
    data[ 8962] = -'sd47592;
    data[ 8963] = -'sd5462;
    data[ 8964] = -'sd38234;
    data[ 8965] =  'sd60044;
    data[ 8966] = -'sd71215;
    data[ 8967] = -'sd6982;
    data[ 8968] = -'sd48874;
    data[ 8969] = -'sd14436;
    data[ 8970] =  'sd62789;
    data[ 8971] = -'sd52000;
    data[ 8972] = -'sd36318;
    data[ 8973] =  'sd73456;
    data[ 8974] =  'sd22669;
    data[ 8975] = -'sd5158;
    data[ 8976] = -'sd36106;
    data[ 8977] =  'sd74940;
    data[ 8978] =  'sd33057;
    data[ 8979] =  'sd67558;
    data[ 8980] = -'sd18617;
    data[ 8981] =  'sd33522;
    data[ 8982] =  'sd70813;
    data[ 8983] =  'sd4168;
    data[ 8984] =  'sd29176;
    data[ 8985] =  'sd40391;
    data[ 8986] = -'sd44945;
    data[ 8987] =  'sd13067;
    data[ 8988] = -'sd72372;
    data[ 8989] = -'sd15081;
    data[ 8990] =  'sd58274;
    data[ 8991] =  'sd80236;
    data[ 8992] =  'sd70129;
    data[ 8993] = -'sd620;
    data[ 8994] = -'sd4340;
    data[ 8995] = -'sd30380;
    data[ 8996] = -'sd48819;
    data[ 8997] = -'sd14051;
    data[ 8998] =  'sd65484;
    data[ 8999] = -'sd33135;
    data[ 9000] = -'sd68104;
    data[ 9001] =  'sd14795;
    data[ 9002] = -'sd60276;
    data[ 9003] =  'sd69591;
    data[ 9004] = -'sd4386;
    data[ 9005] = -'sd30702;
    data[ 9006] = -'sd51073;
    data[ 9007] = -'sd29829;
    data[ 9008] = -'sd44962;
    data[ 9009] =  'sd12948;
    data[ 9010] = -'sd73205;
    data[ 9011] = -'sd20912;
    data[ 9012] =  'sd17457;
    data[ 9013] = -'sd41642;
    data[ 9014] =  'sd36188;
    data[ 9015] = -'sd74366;
    data[ 9016] = -'sd29039;
    data[ 9017] = -'sd39432;
    data[ 9018] =  'sd51658;
    data[ 9019] =  'sd33924;
    data[ 9020] =  'sd73627;
    data[ 9021] =  'sd23866;
    data[ 9022] =  'sd3221;
    data[ 9023] =  'sd22547;
    data[ 9024] = -'sd6012;
    data[ 9025] = -'sd42084;
    data[ 9026] =  'sd33094;
    data[ 9027] =  'sd67817;
    data[ 9028] = -'sd16804;
    data[ 9029] =  'sd46213;
    data[ 9030] = -'sd4191;
    data[ 9031] = -'sd29337;
    data[ 9032] = -'sd41518;
    data[ 9033] =  'sd37056;
    data[ 9034] = -'sd68290;
    data[ 9035] =  'sd13493;
    data[ 9036] = -'sd69390;
    data[ 9037] =  'sd5793;
    data[ 9038] =  'sd40551;
    data[ 9039] = -'sd43825;
    data[ 9040] =  'sd20907;
    data[ 9041] = -'sd17492;
    data[ 9042] =  'sd41397;
    data[ 9043] = -'sd37903;
    data[ 9044] =  'sd62361;
    data[ 9045] = -'sd54996;
    data[ 9046] = -'sd57290;
    data[ 9047] = -'sd73348;
    data[ 9048] = -'sd21913;
    data[ 9049] =  'sd10450;
    data[ 9050] =  'sd73150;
    data[ 9051] =  'sd20527;
    data[ 9052] = -'sd20152;
    data[ 9053] =  'sd22777;
    data[ 9054] = -'sd4402;
    data[ 9055] = -'sd30814;
    data[ 9056] = -'sd51857;
    data[ 9057] = -'sd35317;
    data[ 9058] =  'sd80463;
    data[ 9059] =  'sd71718;
    data[ 9060] =  'sd10503;
    data[ 9061] =  'sd73521;
    data[ 9062] =  'sd23124;
    data[ 9063] = -'sd1973;
    data[ 9064] = -'sd13811;
    data[ 9065] =  'sd67164;
    data[ 9066] = -'sd21375;
    data[ 9067] =  'sd14216;
    data[ 9068] = -'sd64329;
    data[ 9069] =  'sd41220;
    data[ 9070] = -'sd39142;
    data[ 9071] =  'sd53688;
    data[ 9072] =  'sd48134;
    data[ 9073] =  'sd9256;
    data[ 9074] =  'sd64792;
    data[ 9075] = -'sd37979;
    data[ 9076] =  'sd61829;
    data[ 9077] = -'sd58720;
    data[ 9078] =  'sd80483;
    data[ 9079] =  'sd71858;
    data[ 9080] =  'sd11483;
    data[ 9081] =  'sd80381;
    data[ 9082] =  'sd71144;
    data[ 9083] =  'sd6485;
    data[ 9084] =  'sd45395;
    data[ 9085] = -'sd9917;
    data[ 9086] = -'sd69419;
    data[ 9087] =  'sd5590;
    data[ 9088] =  'sd39130;
    data[ 9089] = -'sd53772;
    data[ 9090] = -'sd48722;
    data[ 9091] = -'sd13372;
    data[ 9092] =  'sd70237;
    data[ 9093] =  'sd136;
    data[ 9094] =  'sd952;
    data[ 9095] =  'sd6664;
    data[ 9096] =  'sd46648;
    data[ 9097] = -'sd1146;
    data[ 9098] = -'sd8022;
    data[ 9099] = -'sd56154;
    data[ 9100] = -'sd65396;
    data[ 9101] =  'sd33751;
    data[ 9102] =  'sd72416;
    data[ 9103] =  'sd15389;
    data[ 9104] = -'sd56118;
    data[ 9105] = -'sd65144;
    data[ 9106] =  'sd35515;
    data[ 9107] = -'sd79077;
    data[ 9108] = -'sd62016;
    data[ 9109] =  'sd57411;
    data[ 9110] =  'sd74195;
    data[ 9111] =  'sd27842;
    data[ 9112] =  'sd31053;
    data[ 9113] =  'sd53530;
    data[ 9114] =  'sd47028;
    data[ 9115] =  'sd1514;
    data[ 9116] =  'sd10598;
    data[ 9117] =  'sd74186;
    data[ 9118] =  'sd27779;
    data[ 9119] =  'sd30612;
    data[ 9120] =  'sd50443;
    data[ 9121] =  'sd25419;
    data[ 9122] =  'sd14092;
    data[ 9123] = -'sd65197;
    data[ 9124] =  'sd35144;
    data[ 9125] = -'sd81674;
    data[ 9126] = -'sd80195;
    data[ 9127] = -'sd69842;
    data[ 9128] =  'sd2629;
    data[ 9129] =  'sd18403;
    data[ 9130] = -'sd35020;
    data[ 9131] = -'sd81299;
    data[ 9132] = -'sd77570;
    data[ 9133] = -'sd51467;
    data[ 9134] = -'sd32587;
    data[ 9135] = -'sd64268;
    data[ 9136] =  'sd41647;
    data[ 9137] = -'sd36153;
    data[ 9138] =  'sd74611;
    data[ 9139] =  'sd30754;
    data[ 9140] =  'sd51437;
    data[ 9141] =  'sd32377;
    data[ 9142] =  'sd62798;
    data[ 9143] = -'sd51937;
    data[ 9144] = -'sd35877;
    data[ 9145] =  'sd76543;
    data[ 9146] =  'sd44278;
    data[ 9147] = -'sd17736;
    data[ 9148] =  'sd39689;
    data[ 9149] = -'sd49859;
    data[ 9150] = -'sd21331;
    data[ 9151] =  'sd14524;
    data[ 9152] = -'sd62173;
    data[ 9153] =  'sd56312;
    data[ 9154] =  'sd66502;
    data[ 9155] = -'sd26009;
    data[ 9156] = -'sd18222;
    data[ 9157] =  'sd36287;
    data[ 9158] = -'sd73673;
    data[ 9159] = -'sd24188;
    data[ 9160] = -'sd5475;
    data[ 9161] = -'sd38325;
    data[ 9162] =  'sd59407;
    data[ 9163] = -'sd75674;
    data[ 9164] = -'sd38195;
    data[ 9165] =  'sd60317;
    data[ 9166] = -'sd69304;
    data[ 9167] =  'sd6395;
    data[ 9168] =  'sd44765;
    data[ 9169] = -'sd14327;
    data[ 9170] =  'sd63552;
    data[ 9171] = -'sd46659;
    data[ 9172] =  'sd1069;
    data[ 9173] =  'sd7483;
    data[ 9174] =  'sd52381;
    data[ 9175] =  'sd38985;
    data[ 9176] = -'sd54787;
    data[ 9177] = -'sd55827;
    data[ 9178] = -'sd63107;
    data[ 9179] =  'sd49774;
    data[ 9180] =  'sd20736;
    data[ 9181] = -'sd18689;
    data[ 9182] =  'sd33018;
    data[ 9183] =  'sd67285;
    data[ 9184] = -'sd20528;
    data[ 9185] =  'sd20145;
    data[ 9186] = -'sd22826;
    data[ 9187] =  'sd4059;
    data[ 9188] =  'sd28413;
    data[ 9189] =  'sd35050;
    data[ 9190] =  'sd81509;
    data[ 9191] =  'sd79040;
    data[ 9192] =  'sd61757;
    data[ 9193] = -'sd59224;
    data[ 9194] =  'sd76955;
    data[ 9195] =  'sd47162;
    data[ 9196] =  'sd2452;
    data[ 9197] =  'sd17164;
    data[ 9198] = -'sd43693;
    data[ 9199] =  'sd21831;
    data[ 9200] = -'sd11024;
    data[ 9201] = -'sd77168;
    data[ 9202] = -'sd48653;
    data[ 9203] = -'sd12889;
    data[ 9204] =  'sd73618;
    data[ 9205] =  'sd23803;
    data[ 9206] =  'sd2780;
    data[ 9207] =  'sd19460;
    data[ 9208] = -'sd27621;
    data[ 9209] = -'sd29506;
    data[ 9210] = -'sd42701;
    data[ 9211] =  'sd28775;
    data[ 9212] =  'sd37584;
    data[ 9213] = -'sd64594;
    data[ 9214] =  'sd39365;
    data[ 9215] = -'sd52127;
    data[ 9216] = -'sd37207;
    data[ 9217] =  'sd67233;
    data[ 9218] = -'sd20892;
    data[ 9219] =  'sd17597;
    data[ 9220] = -'sd40662;
    data[ 9221] =  'sd43048;
    data[ 9222] = -'sd26346;
    data[ 9223] = -'sd20581;
    data[ 9224] =  'sd19774;
    data[ 9225] = -'sd25423;
    data[ 9226] = -'sd14120;
    data[ 9227] =  'sd65001;
    data[ 9228] = -'sd36516;
    data[ 9229] =  'sd72070;
    data[ 9230] =  'sd12967;
    data[ 9231] = -'sd73072;
    data[ 9232] = -'sd19981;
    data[ 9233] =  'sd23974;
    data[ 9234] =  'sd3977;
    data[ 9235] =  'sd27839;
    data[ 9236] =  'sd31032;
    data[ 9237] =  'sd53383;
    data[ 9238] =  'sd45999;
    data[ 9239] = -'sd5689;
    data[ 9240] = -'sd39823;
    data[ 9241] =  'sd48921;
    data[ 9242] =  'sd14765;
    data[ 9243] = -'sd60486;
    data[ 9244] =  'sd68121;
    data[ 9245] = -'sd14676;
    data[ 9246] =  'sd61109;
    data[ 9247] = -'sd63760;
    data[ 9248] =  'sd45203;
    data[ 9249] = -'sd11261;
    data[ 9250] = -'sd78827;
    data[ 9251] = -'sd60266;
    data[ 9252] =  'sd69661;
    data[ 9253] = -'sd3896;
    data[ 9254] = -'sd27272;
    data[ 9255] = -'sd27063;
    data[ 9256] = -'sd25600;
    data[ 9257] = -'sd15359;
    data[ 9258] =  'sd56328;
    data[ 9259] =  'sd66614;
    data[ 9260] = -'sd25225;
    data[ 9261] = -'sd12734;
    data[ 9262] =  'sd74703;
    data[ 9263] =  'sd31398;
    data[ 9264] =  'sd55945;
    data[ 9265] =  'sd63933;
    data[ 9266] = -'sd43992;
    data[ 9267] =  'sd19738;
    data[ 9268] = -'sd25675;
    data[ 9269] = -'sd15884;
    data[ 9270] =  'sd52653;
    data[ 9271] =  'sd40889;
    data[ 9272] = -'sd41459;
    data[ 9273] =  'sd37469;
    data[ 9274] = -'sd65399;
    data[ 9275] =  'sd33730;
    data[ 9276] =  'sd72269;
    data[ 9277] =  'sd14360;
    data[ 9278] = -'sd63321;
    data[ 9279] =  'sd48276;
    data[ 9280] =  'sd10250;
    data[ 9281] =  'sd71750;
    data[ 9282] =  'sd10727;
    data[ 9283] =  'sd75089;
    data[ 9284] =  'sd34100;
    data[ 9285] =  'sd74859;
    data[ 9286] =  'sd32490;
    data[ 9287] =  'sd63589;
    data[ 9288] = -'sd46400;
    data[ 9289] =  'sd2882;
    data[ 9290] =  'sd20174;
    data[ 9291] = -'sd22623;
    data[ 9292] =  'sd5480;
    data[ 9293] =  'sd38360;
    data[ 9294] = -'sd59162;
    data[ 9295] =  'sd77389;
    data[ 9296] =  'sd50200;
    data[ 9297] =  'sd23718;
    data[ 9298] =  'sd2185;
    data[ 9299] =  'sd15295;
    data[ 9300] = -'sd56776;
    data[ 9301] = -'sd69750;
    data[ 9302] =  'sd3273;
    data[ 9303] =  'sd22911;
    data[ 9304] = -'sd3464;
    data[ 9305] = -'sd24248;
    data[ 9306] = -'sd5895;
    data[ 9307] = -'sd41265;
    data[ 9308] =  'sd38827;
    data[ 9309] = -'sd55893;
    data[ 9310] = -'sd63569;
    data[ 9311] =  'sd46540;
    data[ 9312] = -'sd1902;
    data[ 9313] = -'sd13314;
    data[ 9314] =  'sd70643;
    data[ 9315] =  'sd2978;
    data[ 9316] =  'sd20846;
    data[ 9317] = -'sd17919;
    data[ 9318] =  'sd38408;
    data[ 9319] = -'sd58826;
    data[ 9320] =  'sd79741;
    data[ 9321] =  'sd66664;
    data[ 9322] = -'sd24875;
    data[ 9323] = -'sd10284;
    data[ 9324] = -'sd71988;
    data[ 9325] = -'sd12393;
    data[ 9326] =  'sd77090;
    data[ 9327] =  'sd48107;
    data[ 9328] =  'sd9067;
    data[ 9329] =  'sd63469;
    data[ 9330] = -'sd47240;
    data[ 9331] = -'sd2998;
    data[ 9332] = -'sd20986;
    data[ 9333] =  'sd16939;
    data[ 9334] = -'sd45268;
    data[ 9335] =  'sd10806;
    data[ 9336] =  'sd75642;
    data[ 9337] =  'sd37971;
    data[ 9338] = -'sd61885;
    data[ 9339] =  'sd58328;
    data[ 9340] =  'sd80614;
    data[ 9341] =  'sd72775;
    data[ 9342] =  'sd17902;
    data[ 9343] = -'sd38527;
    data[ 9344] =  'sd57993;
    data[ 9345] =  'sd78269;
    data[ 9346] =  'sd56360;
    data[ 9347] =  'sd66838;
    data[ 9348] = -'sd23657;
    data[ 9349] = -'sd1758;
    data[ 9350] = -'sd12306;
    data[ 9351] =  'sd77699;
    data[ 9352] =  'sd52370;
    data[ 9353] =  'sd38908;
    data[ 9354] = -'sd55326;
    data[ 9355] = -'sd59600;
    data[ 9356] =  'sd74323;
    data[ 9357] =  'sd28738;
    data[ 9358] =  'sd37325;
    data[ 9359] = -'sd66407;
    data[ 9360] =  'sd26674;
    data[ 9361] =  'sd22877;
    data[ 9362] = -'sd3702;
    data[ 9363] = -'sd25914;
    data[ 9364] = -'sd17557;
    data[ 9365] =  'sd40942;
    data[ 9366] = -'sd41088;
    data[ 9367] =  'sd40066;
    data[ 9368] = -'sd47220;
    data[ 9369] = -'sd2858;
    data[ 9370] = -'sd20006;
    data[ 9371] =  'sd23799;
    data[ 9372] =  'sd2752;
    data[ 9373] =  'sd19264;
    data[ 9374] = -'sd28993;
    data[ 9375] = -'sd39110;
    data[ 9376] =  'sd53912;
    data[ 9377] =  'sd49702;
    data[ 9378] =  'sd20232;
    data[ 9379] = -'sd22217;
    data[ 9380] =  'sd8322;
    data[ 9381] =  'sd58254;
    data[ 9382] =  'sd80096;
    data[ 9383] =  'sd69149;
    data[ 9384] = -'sd7480;
    data[ 9385] = -'sd52360;
    data[ 9386] = -'sd38838;
    data[ 9387] =  'sd55816;
    data[ 9388] =  'sd63030;
    data[ 9389] = -'sd50313;
    data[ 9390] = -'sd24509;
    data[ 9391] = -'sd7722;
    data[ 9392] = -'sd54054;
    data[ 9393] = -'sd50696;
    data[ 9394] = -'sd27190;
    data[ 9395] = -'sd26489;
    data[ 9396] = -'sd21582;
    data[ 9397] =  'sd12767;
    data[ 9398] = -'sd74472;
    data[ 9399] = -'sd29781;
    data[ 9400] = -'sd44626;
    data[ 9401] =  'sd15300;
    data[ 9402] = -'sd56741;
    data[ 9403] = -'sd69505;
    data[ 9404] =  'sd4988;
    data[ 9405] =  'sd34916;
    data[ 9406] =  'sd80571;
    data[ 9407] =  'sd72474;
    data[ 9408] =  'sd15795;
    data[ 9409] = -'sd53276;
    data[ 9410] = -'sd45250;
    data[ 9411] =  'sd10932;
    data[ 9412] =  'sd76524;
    data[ 9413] =  'sd44145;
    data[ 9414] = -'sd18667;
    data[ 9415] =  'sd33172;
    data[ 9416] =  'sd68363;
    data[ 9417] = -'sd12982;
    data[ 9418] =  'sd72967;
    data[ 9419] =  'sd19246;
    data[ 9420] = -'sd29119;
    data[ 9421] = -'sd39992;
    data[ 9422] =  'sd47738;
    data[ 9423] =  'sd6484;
    data[ 9424] =  'sd45388;
    data[ 9425] = -'sd9966;
    data[ 9426] = -'sd69762;
    data[ 9427] =  'sd3189;
    data[ 9428] =  'sd22323;
    data[ 9429] = -'sd7580;
    data[ 9430] = -'sd53060;
    data[ 9431] = -'sd43738;
    data[ 9432] =  'sd21516;
    data[ 9433] = -'sd13229;
    data[ 9434] =  'sd71238;
    data[ 9435] =  'sd7143;
    data[ 9436] =  'sd50001;
    data[ 9437] =  'sd22325;
    data[ 9438] = -'sd7566;
    data[ 9439] = -'sd52962;
    data[ 9440] = -'sd43052;
    data[ 9441] =  'sd26318;
    data[ 9442] =  'sd20385;
    data[ 9443] = -'sd21146;
    data[ 9444] =  'sd15819;
    data[ 9445] = -'sd53108;
    data[ 9446] = -'sd44074;
    data[ 9447] =  'sd19164;
    data[ 9448] = -'sd29693;
    data[ 9449] = -'sd44010;
    data[ 9450] =  'sd19612;
    data[ 9451] = -'sd26557;
    data[ 9452] = -'sd22058;
    data[ 9453] =  'sd9435;
    data[ 9454] =  'sd66045;
    data[ 9455] = -'sd29208;
    data[ 9456] = -'sd40615;
    data[ 9457] =  'sd43377;
    data[ 9458] = -'sd24043;
    data[ 9459] = -'sd4460;
    data[ 9460] = -'sd31220;
    data[ 9461] = -'sd54699;
    data[ 9462] = -'sd55211;
    data[ 9463] = -'sd58795;
    data[ 9464] =  'sd79958;
    data[ 9465] =  'sd68183;
    data[ 9466] = -'sd14242;
    data[ 9467] =  'sd64147;
    data[ 9468] = -'sd42494;
    data[ 9469] =  'sd30224;
    data[ 9470] =  'sd47727;
    data[ 9471] =  'sd6407;
    data[ 9472] =  'sd44849;
    data[ 9473] = -'sd13739;
    data[ 9474] =  'sd67668;
    data[ 9475] = -'sd17847;
    data[ 9476] =  'sd38912;
    data[ 9477] = -'sd55298;
    data[ 9478] = -'sd59404;
    data[ 9479] =  'sd75695;
    data[ 9480] =  'sd38342;
    data[ 9481] = -'sd59288;
    data[ 9482] =  'sd76507;
    data[ 9483] =  'sd44026;
    data[ 9484] = -'sd19500;
    data[ 9485] =  'sd27341;
    data[ 9486] =  'sd27546;
    data[ 9487] =  'sd28981;
    data[ 9488] =  'sd39026;
    data[ 9489] = -'sd54500;
    data[ 9490] = -'sd53818;
    data[ 9491] = -'sd49044;
    data[ 9492] = -'sd15626;
    data[ 9493] =  'sd54459;
    data[ 9494] =  'sd53531;
    data[ 9495] =  'sd47035;
    data[ 9496] =  'sd1563;
    data[ 9497] =  'sd10941;
    data[ 9498] =  'sd76587;
    data[ 9499] =  'sd44586;
    data[ 9500] = -'sd15580;
    data[ 9501] =  'sd54781;
    data[ 9502] =  'sd55785;
    data[ 9503] =  'sd62813;
    data[ 9504] = -'sd51832;
    data[ 9505] = -'sd35142;
    data[ 9506] =  'sd81688;
    data[ 9507] =  'sd80293;
    data[ 9508] =  'sd70528;
    data[ 9509] =  'sd2173;
    data[ 9510] =  'sd15211;
    data[ 9511] = -'sd57364;
    data[ 9512] = -'sd73866;
    data[ 9513] = -'sd25539;
    data[ 9514] = -'sd14932;
    data[ 9515] =  'sd59317;
    data[ 9516] = -'sd76304;
    data[ 9517] = -'sd42605;
    data[ 9518] =  'sd29447;
    data[ 9519] =  'sd42288;
    data[ 9520] = -'sd31666;
    data[ 9521] = -'sd57821;
    data[ 9522] = -'sd77065;
    data[ 9523] = -'sd47932;
    data[ 9524] = -'sd7842;
    data[ 9525] = -'sd54894;
    data[ 9526] = -'sd56576;
    data[ 9527] = -'sd68350;
    data[ 9528] =  'sd13073;
    data[ 9529] = -'sd72330;
    data[ 9530] = -'sd14787;
    data[ 9531] =  'sd60332;
    data[ 9532] = -'sd69199;
    data[ 9533] =  'sd7130;
    data[ 9534] =  'sd49910;
    data[ 9535] =  'sd21688;
    data[ 9536] = -'sd12025;
    data[ 9537] =  'sd79666;
    data[ 9538] =  'sd66139;
    data[ 9539] = -'sd28550;
    data[ 9540] = -'sd36009;
    data[ 9541] =  'sd75619;
    data[ 9542] =  'sd37810;
    data[ 9543] = -'sd63012;
    data[ 9544] =  'sd50439;
    data[ 9545] =  'sd25391;
    data[ 9546] =  'sd13896;
    data[ 9547] = -'sd66569;
    data[ 9548] =  'sd25540;
    data[ 9549] =  'sd14939;
    data[ 9550] = -'sd59268;
    data[ 9551] =  'sd76647;
    data[ 9552] =  'sd45006;
    data[ 9553] = -'sd12640;
    data[ 9554] =  'sd75361;
    data[ 9555] =  'sd36004;
    data[ 9556] = -'sd75654;
    data[ 9557] = -'sd38055;
    data[ 9558] =  'sd61297;
    data[ 9559] = -'sd62444;
    data[ 9560] =  'sd54415;
    data[ 9561] =  'sd53223;
    data[ 9562] =  'sd44879;
    data[ 9563] = -'sd13529;
    data[ 9564] =  'sd69138;
    data[ 9565] = -'sd7557;
    data[ 9566] = -'sd52899;
    data[ 9567] = -'sd42611;
    data[ 9568] =  'sd29405;
    data[ 9569] =  'sd41994;
    data[ 9570] = -'sd33724;
    data[ 9571] = -'sd72227;
    data[ 9572] = -'sd14066;
    data[ 9573] =  'sd65379;
    data[ 9574] = -'sd33870;
    data[ 9575] = -'sd73249;
    data[ 9576] = -'sd21220;
    data[ 9577] =  'sd15301;
    data[ 9578] = -'sd56734;
    data[ 9579] = -'sd69456;
    data[ 9580] =  'sd5331;
    data[ 9581] =  'sd37317;
    data[ 9582] = -'sd66463;
    data[ 9583] =  'sd26282;
    data[ 9584] =  'sd20133;
    data[ 9585] = -'sd22910;
    data[ 9586] =  'sd3471;
    data[ 9587] =  'sd24297;
    data[ 9588] =  'sd6238;
    data[ 9589] =  'sd43666;
    data[ 9590] = -'sd22020;
    data[ 9591] =  'sd9701;
    data[ 9592] =  'sd67907;
    data[ 9593] = -'sd16174;
    data[ 9594] =  'sd50623;
    data[ 9595] =  'sd26679;
    data[ 9596] =  'sd22912;
    data[ 9597] = -'sd3457;
    data[ 9598] = -'sd24199;
    data[ 9599] = -'sd5552;
    data[ 9600] = -'sd38864;
    data[ 9601] =  'sd55634;
    data[ 9602] =  'sd61756;
    data[ 9603] = -'sd59231;
    data[ 9604] =  'sd76906;
    data[ 9605] =  'sd46819;
    data[ 9606] =  'sd51;
    data[ 9607] =  'sd357;
    data[ 9608] =  'sd2499;
    data[ 9609] =  'sd17493;
    data[ 9610] = -'sd41390;
    data[ 9611] =  'sd37952;
    data[ 9612] = -'sd62018;
    data[ 9613] =  'sd57397;
    data[ 9614] =  'sd74097;
    data[ 9615] =  'sd27156;
    data[ 9616] =  'sd26251;
    data[ 9617] =  'sd19916;
    data[ 9618] = -'sd24429;
    data[ 9619] = -'sd7162;
    data[ 9620] = -'sd50134;
    data[ 9621] = -'sd23256;
    data[ 9622] =  'sd1049;
    data[ 9623] =  'sd7343;
    data[ 9624] =  'sd51401;
    data[ 9625] =  'sd32125;
    data[ 9626] =  'sd61034;
    data[ 9627] = -'sd64285;
    data[ 9628] =  'sd41528;
    data[ 9629] = -'sd36986;
    data[ 9630] =  'sd68780;
    data[ 9631] = -'sd10063;
    data[ 9632] = -'sd70441;
    data[ 9633] = -'sd1564;
    data[ 9634] = -'sd10948;
    data[ 9635] = -'sd76636;
    data[ 9636] = -'sd44929;
    data[ 9637] =  'sd13179;
    data[ 9638] = -'sd71588;
    data[ 9639] = -'sd9593;
    data[ 9640] = -'sd67151;
    data[ 9641] =  'sd21466;
    data[ 9642] = -'sd13579;
    data[ 9643] =  'sd68788;
    data[ 9644] = -'sd10007;
    data[ 9645] = -'sd70049;
    data[ 9646] =  'sd1180;
    data[ 9647] =  'sd8260;
    data[ 9648] =  'sd57820;
    data[ 9649] =  'sd77058;
    data[ 9650] =  'sd47883;
    data[ 9651] =  'sd7499;
    data[ 9652] =  'sd52493;
    data[ 9653] =  'sd39769;
    data[ 9654] = -'sd49299;
    data[ 9655] = -'sd17411;
    data[ 9656] =  'sd41964;
    data[ 9657] = -'sd33934;
    data[ 9658] = -'sd73697;
    data[ 9659] = -'sd24356;
    data[ 9660] = -'sd6651;
    data[ 9661] = -'sd46557;
    data[ 9662] =  'sd1783;
    data[ 9663] =  'sd12481;
    data[ 9664] = -'sd76474;
    data[ 9665] = -'sd43795;
    data[ 9666] =  'sd21117;
    data[ 9667] = -'sd16022;
    data[ 9668] =  'sd51687;
    data[ 9669] =  'sd34127;
    data[ 9670] =  'sd75048;
    data[ 9671] =  'sd33813;
    data[ 9672] =  'sd72850;
    data[ 9673] =  'sd18427;
    data[ 9674] = -'sd34852;
    data[ 9675] = -'sd80123;
    data[ 9676] = -'sd69338;
    data[ 9677] =  'sd6157;
    data[ 9678] =  'sd43099;
    data[ 9679] = -'sd25989;
    data[ 9680] = -'sd18082;
    data[ 9681] =  'sd37267;
    data[ 9682] = -'sd66813;
    data[ 9683] =  'sd23832;
    data[ 9684] =  'sd2983;
    data[ 9685] =  'sd20881;
    data[ 9686] = -'sd17674;
    data[ 9687] =  'sd40123;
    data[ 9688] = -'sd46821;
    data[ 9689] = -'sd65;
    data[ 9690] = -'sd455;
    data[ 9691] = -'sd3185;
    data[ 9692] = -'sd22295;
    data[ 9693] =  'sd7776;
    data[ 9694] =  'sd54432;
    data[ 9695] =  'sd53342;
    data[ 9696] =  'sd45712;
    data[ 9697] = -'sd7698;
    data[ 9698] = -'sd53886;
    data[ 9699] = -'sd49520;
    data[ 9700] = -'sd18958;
    data[ 9701] =  'sd31135;
    data[ 9702] =  'sd54104;
    data[ 9703] =  'sd51046;
    data[ 9704] =  'sd29640;
    data[ 9705] =  'sd43639;
    data[ 9706] = -'sd22209;
    data[ 9707] =  'sd8378;
    data[ 9708] =  'sd58646;
    data[ 9709] = -'sd81001;
    data[ 9710] = -'sd75484;
    data[ 9711] = -'sd36865;
    data[ 9712] =  'sd69627;
    data[ 9713] = -'sd4134;
    data[ 9714] = -'sd28938;
    data[ 9715] = -'sd38725;
    data[ 9716] =  'sd56607;
    data[ 9717] =  'sd68567;
    data[ 9718] = -'sd11554;
    data[ 9719] = -'sd80878;
    data[ 9720] = -'sd74623;
    data[ 9721] = -'sd30838;
    data[ 9722] = -'sd52025;
    data[ 9723] = -'sd36493;
    data[ 9724] =  'sd72231;
    data[ 9725] =  'sd14094;
    data[ 9726] = -'sd65183;
    data[ 9727] =  'sd35242;
    data[ 9728] = -'sd80988;
    data[ 9729] = -'sd75393;
    data[ 9730] = -'sd36228;
    data[ 9731] =  'sd74086;
    data[ 9732] =  'sd27079;
    data[ 9733] =  'sd25712;
    data[ 9734] =  'sd16143;
    data[ 9735] = -'sd50840;
    data[ 9736] = -'sd28198;
    data[ 9737] = -'sd33545;
    data[ 9738] = -'sd70974;
    data[ 9739] = -'sd5295;
    data[ 9740] = -'sd37065;
    data[ 9741] =  'sd68227;
    data[ 9742] = -'sd13934;
    data[ 9743] =  'sd66303;
    data[ 9744] = -'sd27402;
    data[ 9745] = -'sd27973;
    data[ 9746] = -'sd31970;
    data[ 9747] = -'sd59949;
    data[ 9748] =  'sd71880;
    data[ 9749] =  'sd11637;
    data[ 9750] =  'sd81459;
    data[ 9751] =  'sd78690;
    data[ 9752] =  'sd59307;
    data[ 9753] = -'sd76374;
    data[ 9754] = -'sd43095;
    data[ 9755] =  'sd26017;
    data[ 9756] =  'sd18278;
    data[ 9757] = -'sd35895;
    data[ 9758] =  'sd76417;
    data[ 9759] =  'sd43396;
    data[ 9760] = -'sd23910;
    data[ 9761] = -'sd3529;
    data[ 9762] = -'sd24703;
    data[ 9763] = -'sd9080;
    data[ 9764] = -'sd63560;
    data[ 9765] =  'sd46603;
    data[ 9766] = -'sd1461;
    data[ 9767] = -'sd10227;
    data[ 9768] = -'sd71589;
    data[ 9769] = -'sd9600;
    data[ 9770] = -'sd67200;
    data[ 9771] =  'sd21123;
    data[ 9772] = -'sd15980;
    data[ 9773] =  'sd51981;
    data[ 9774] =  'sd36185;
    data[ 9775] = -'sd74387;
    data[ 9776] = -'sd29186;
    data[ 9777] = -'sd40461;
    data[ 9778] =  'sd44455;
    data[ 9779] = -'sd16497;
    data[ 9780] =  'sd48362;
    data[ 9781] =  'sd10852;
    data[ 9782] =  'sd75964;
    data[ 9783] =  'sd40225;
    data[ 9784] = -'sd46107;
    data[ 9785] =  'sd4933;
    data[ 9786] =  'sd34531;
    data[ 9787] =  'sd77876;
    data[ 9788] =  'sd53609;
    data[ 9789] =  'sd47581;
    data[ 9790] =  'sd5385;
    data[ 9791] =  'sd37695;
    data[ 9792] = -'sd63817;
    data[ 9793] =  'sd44804;
    data[ 9794] = -'sd14054;
    data[ 9795] =  'sd65463;
    data[ 9796] = -'sd33282;
    data[ 9797] = -'sd69133;
    data[ 9798] =  'sd7592;
    data[ 9799] =  'sd53144;
    data[ 9800] =  'sd44326;
    data[ 9801] = -'sd17400;
    data[ 9802] =  'sd42041;
    data[ 9803] = -'sd33395;
    data[ 9804] = -'sd69924;
    data[ 9805] =  'sd2055;
    data[ 9806] =  'sd14385;
    data[ 9807] = -'sd63146;
    data[ 9808] =  'sd49501;
    data[ 9809] =  'sd18825;
    data[ 9810] = -'sd32066;
    data[ 9811] = -'sd60621;
    data[ 9812] =  'sd67176;
    data[ 9813] = -'sd21291;
    data[ 9814] =  'sd14804;
    data[ 9815] = -'sd60213;
    data[ 9816] =  'sd70032;
    data[ 9817] = -'sd1299;
    data[ 9818] = -'sd9093;
    data[ 9819] = -'sd63651;
    data[ 9820] =  'sd45966;
    data[ 9821] = -'sd5920;
    data[ 9822] = -'sd41440;
    data[ 9823] =  'sd37602;
    data[ 9824] = -'sd64468;
    data[ 9825] =  'sd40247;
    data[ 9826] = -'sd45953;
    data[ 9827] =  'sd6011;
    data[ 9828] =  'sd42077;
    data[ 9829] = -'sd33143;
    data[ 9830] = -'sd68160;
    data[ 9831] =  'sd14403;
    data[ 9832] = -'sd63020;
    data[ 9833] =  'sd50383;
    data[ 9834] =  'sd24999;
    data[ 9835] =  'sd11152;
    data[ 9836] =  'sd78064;
    data[ 9837] =  'sd54925;
    data[ 9838] =  'sd56793;
    data[ 9839] =  'sd69869;
    data[ 9840] = -'sd2440;
    data[ 9841] = -'sd17080;
    data[ 9842] =  'sd44281;
    data[ 9843] = -'sd17715;
    data[ 9844] =  'sd39836;
    data[ 9845] = -'sd48830;
    data[ 9846] = -'sd14128;
    data[ 9847] =  'sd64945;
    data[ 9848] = -'sd36908;
    data[ 9849] =  'sd69326;
    data[ 9850] = -'sd6241;
    data[ 9851] = -'sd43687;
    data[ 9852] =  'sd21873;
    data[ 9853] = -'sd10730;
    data[ 9854] = -'sd75110;
    data[ 9855] = -'sd34247;
    data[ 9856] = -'sd75888;
    data[ 9857] = -'sd39693;
    data[ 9858] =  'sd49831;
    data[ 9859] =  'sd21135;
    data[ 9860] = -'sd15896;
    data[ 9861] =  'sd52569;
    data[ 9862] =  'sd40301;
    data[ 9863] = -'sd45575;
    data[ 9864] =  'sd8657;
    data[ 9865] =  'sd60599;
    data[ 9866] = -'sd67330;
    data[ 9867] =  'sd20213;
    data[ 9868] = -'sd22350;
    data[ 9869] =  'sd7391;
    data[ 9870] =  'sd51737;
    data[ 9871] =  'sd34477;
    data[ 9872] =  'sd77498;
    data[ 9873] =  'sd50963;
    data[ 9874] =  'sd29059;
    data[ 9875] =  'sd39572;
    data[ 9876] = -'sd50678;
    data[ 9877] = -'sd27064;
    data[ 9878] = -'sd25607;
    data[ 9879] = -'sd15408;
    data[ 9880] =  'sd55985;
    data[ 9881] =  'sd64213;
    data[ 9882] = -'sd42032;
    data[ 9883] =  'sd33458;
    data[ 9884] =  'sd70365;
    data[ 9885] =  'sd1032;
    data[ 9886] =  'sd7224;
    data[ 9887] =  'sd50568;
    data[ 9888] =  'sd26294;
    data[ 9889] =  'sd20217;
    data[ 9890] = -'sd22322;
    data[ 9891] =  'sd7587;
    data[ 9892] =  'sd53109;
    data[ 9893] =  'sd44081;
    data[ 9894] = -'sd19115;
    data[ 9895] =  'sd30036;
    data[ 9896] =  'sd46411;
    data[ 9897] = -'sd2805;
    data[ 9898] = -'sd19635;
    data[ 9899] =  'sd26396;
    data[ 9900] =  'sd20931;
    data[ 9901] = -'sd17324;
    data[ 9902] =  'sd42573;
    data[ 9903] = -'sd29671;
    data[ 9904] = -'sd43856;
    data[ 9905] =  'sd20690;
    data[ 9906] = -'sd19011;
    data[ 9907] =  'sd30764;
    data[ 9908] =  'sd51507;
    data[ 9909] =  'sd32867;
    data[ 9910] =  'sd66228;
    data[ 9911] = -'sd27927;
    data[ 9912] = -'sd31648;
    data[ 9913] = -'sd57695;
    data[ 9914] = -'sd76183;
    data[ 9915] = -'sd41758;
    data[ 9916] =  'sd35376;
    data[ 9917] = -'sd80050;
    data[ 9918] = -'sd68827;
    data[ 9919] =  'sd9734;
    data[ 9920] =  'sd68138;
    data[ 9921] = -'sd14557;
    data[ 9922] =  'sd61942;
    data[ 9923] = -'sd57929;
    data[ 9924] = -'sd77821;
    data[ 9925] = -'sd53224;
    data[ 9926] = -'sd44886;
    data[ 9927] =  'sd13480;
    data[ 9928] = -'sd69481;
    data[ 9929] =  'sd5156;
    data[ 9930] =  'sd36092;
    data[ 9931] = -'sd75038;
    data[ 9932] = -'sd33743;
    data[ 9933] = -'sd72360;
    data[ 9934] = -'sd14997;
    data[ 9935] =  'sd58862;
    data[ 9936] = -'sd79489;
    data[ 9937] = -'sd64900;
    data[ 9938] =  'sd37223;
    data[ 9939] = -'sd67121;
    data[ 9940] =  'sd21676;
    data[ 9941] = -'sd12109;
    data[ 9942] =  'sd79078;
    data[ 9943] =  'sd62023;
    data[ 9944] = -'sd57362;
    data[ 9945] = -'sd73852;
    data[ 9946] = -'sd25441;
    data[ 9947] = -'sd14246;
    data[ 9948] =  'sd64119;
    data[ 9949] = -'sd42690;
    data[ 9950] =  'sd28852;
    data[ 9951] =  'sd38123;
    data[ 9952] = -'sd60821;
    data[ 9953] =  'sd65776;
    data[ 9954] = -'sd31091;
    data[ 9955] = -'sd53796;
    data[ 9956] = -'sd48890;
    data[ 9957] = -'sd14548;
    data[ 9958] =  'sd62005;
    data[ 9959] = -'sd57488;
    data[ 9960] = -'sd74734;
    data[ 9961] = -'sd31615;
    data[ 9962] = -'sd57464;
    data[ 9963] = -'sd74566;
    data[ 9964] = -'sd30439;
    data[ 9965] = -'sd49232;
    data[ 9966] = -'sd16942;
    data[ 9967] =  'sd45247;
    data[ 9968] = -'sd10953;
    data[ 9969] = -'sd76671;
    data[ 9970] = -'sd45174;
    data[ 9971] =  'sd11464;
    data[ 9972] =  'sd80248;
    data[ 9973] =  'sd70213;
    data[ 9974] = -'sd32;
    data[ 9975] = -'sd224;
    data[ 9976] = -'sd1568;
    data[ 9977] = -'sd10976;
    data[ 9978] = -'sd76832;
    data[ 9979] = -'sd46301;
    data[ 9980] =  'sd3575;
    data[ 9981] =  'sd25025;
    data[ 9982] =  'sd11334;
    data[ 9983] =  'sd79338;
    data[ 9984] =  'sd63843;
    data[ 9985] = -'sd44622;
    data[ 9986] =  'sd15328;
    data[ 9987] = -'sd56545;
    data[ 9988] = -'sd68133;
    data[ 9989] =  'sd14592;
    data[ 9990] = -'sd61697;
    data[ 9991] =  'sd59644;
    data[ 9992] = -'sd74015;
    data[ 9993] = -'sd26582;
    data[ 9994] = -'sd22233;
    data[ 9995] =  'sd8210;
    data[ 9996] =  'sd57470;
    data[ 9997] =  'sd74608;
    data[ 9998] =  'sd30733;
    data[ 9999] =  'sd51290;
    data[10000] =  'sd31348;
    data[10001] =  'sd55595;
    data[10002] =  'sd61483;
    data[10003] = -'sd61142;
    data[10004] =  'sd63529;
    data[10005] = -'sd46820;
    data[10006] = -'sd58;
    data[10007] = -'sd406;
    data[10008] = -'sd2842;
    data[10009] = -'sd19894;
    data[10010] =  'sd24583;
    data[10011] =  'sd8240;
    data[10012] =  'sd57680;
    data[10013] =  'sd76078;
    data[10014] =  'sd41023;
    data[10015] = -'sd40521;
    data[10016] =  'sd44035;
    data[10017] = -'sd19437;
    data[10018] =  'sd27782;
    data[10019] =  'sd30633;
    data[10020] =  'sd50590;
    data[10021] =  'sd26448;
    data[10022] =  'sd21295;
    data[10023] = -'sd14776;
    data[10024] =  'sd60409;
    data[10025] = -'sd68660;
    data[10026] =  'sd10903;
    data[10027] =  'sd76321;
    data[10028] =  'sd42724;
    data[10029] = -'sd28614;
    data[10030] = -'sd36457;
    data[10031] =  'sd72483;
    data[10032] =  'sd15858;
    data[10033] = -'sd52835;
    data[10034] = -'sd42163;
    data[10035] =  'sd32541;
    data[10036] =  'sd63946;
    data[10037] = -'sd43901;
    data[10038] =  'sd20375;
    data[10039] = -'sd21216;
    data[10040] =  'sd15329;
    data[10041] = -'sd56538;
    data[10042] = -'sd68084;
    data[10043] =  'sd14935;
    data[10044] = -'sd59296;
    data[10045] =  'sd76451;
    data[10046] =  'sd43634;
    data[10047] = -'sd22244;
    data[10048] =  'sd8133;
    data[10049] =  'sd56931;
    data[10050] =  'sd70835;
    data[10051] =  'sd4322;
    data[10052] =  'sd30254;
    data[10053] =  'sd47937;
    data[10054] =  'sd7877;
    data[10055] =  'sd55139;
    data[10056] =  'sd58291;
    data[10057] =  'sd80355;
    data[10058] =  'sd70962;
    data[10059] =  'sd5211;
    data[10060] =  'sd36477;
    data[10061] = -'sd72343;
    data[10062] = -'sd14878;
    data[10063] =  'sd59695;
    data[10064] = -'sd73658;
    data[10065] = -'sd24083;
    data[10066] = -'sd4740;
    data[10067] = -'sd33180;
    data[10068] = -'sd68419;
    data[10069] =  'sd12590;
    data[10070] = -'sd75711;
    data[10071] = -'sd38454;
    data[10072] =  'sd58504;
    data[10073] =  'sd81846;
    data[10074] =  'sd81399;
    data[10075] =  'sd78270;
    data[10076] =  'sd56367;
    data[10077] =  'sd66887;
    data[10078] = -'sd23314;
    data[10079] =  'sd643;
    data[10080] =  'sd4501;
    data[10081] =  'sd31507;
    data[10082] =  'sd56708;
    data[10083] =  'sd69274;
    data[10084] = -'sd6605;
    data[10085] = -'sd46235;
    data[10086] =  'sd4037;
    data[10087] =  'sd28259;
    data[10088] =  'sd33972;
    data[10089] =  'sd73963;
    data[10090] =  'sd26218;
    data[10091] =  'sd19685;
    data[10092] = -'sd26046;
    data[10093] = -'sd18481;
    data[10094] =  'sd34474;
    data[10095] =  'sd77477;
    data[10096] =  'sd50816;
    data[10097] =  'sd28030;
    data[10098] =  'sd32369;
    data[10099] =  'sd62742;
    data[10100] = -'sd52329;
    data[10101] = -'sd38621;
    data[10102] =  'sd57335;
    data[10103] =  'sd73663;
    data[10104] =  'sd24118;
    data[10105] =  'sd4985;
    data[10106] =  'sd34895;
    data[10107] =  'sd80424;
    data[10108] =  'sd71445;
    data[10109] =  'sd8592;
    data[10110] =  'sd60144;
    data[10111] = -'sd70515;
    data[10112] = -'sd2082;
    data[10113] = -'sd14574;
    data[10114] =  'sd61823;
    data[10115] = -'sd58762;
    data[10116] =  'sd80189;
    data[10117] =  'sd69800;
    data[10118] = -'sd2923;
    data[10119] = -'sd20461;
    data[10120] =  'sd20614;
    data[10121] = -'sd19543;
    data[10122] =  'sd27040;
    data[10123] =  'sd25439;
    data[10124] =  'sd14232;
    data[10125] = -'sd64217;
    data[10126] =  'sd42004;
    data[10127] = -'sd33654;
    data[10128] = -'sd71737;
    data[10129] = -'sd10636;
    data[10130] = -'sd74452;
    data[10131] = -'sd29641;
    data[10132] = -'sd43646;
    data[10133] =  'sd22160;
    data[10134] = -'sd8721;
    data[10135] = -'sd61047;
    data[10136] =  'sd64194;
    data[10137] = -'sd42165;
    data[10138] =  'sd32527;
    data[10139] =  'sd63848;
    data[10140] = -'sd44587;
    data[10141] =  'sd15573;
    data[10142] = -'sd54830;
    data[10143] = -'sd56128;
    data[10144] = -'sd65214;
    data[10145] =  'sd35025;
    data[10146] =  'sd81334;
    data[10147] =  'sd77815;
    data[10148] =  'sd53182;
    data[10149] =  'sd44592;
    data[10150] = -'sd15538;
    data[10151] =  'sd55075;
    data[10152] =  'sd57843;
    data[10153] =  'sd77219;
    data[10154] =  'sd49010;
    data[10155] =  'sd15388;
    data[10156] = -'sd56125;
    data[10157] = -'sd65193;
    data[10158] =  'sd35172;
    data[10159] = -'sd81478;
    data[10160] = -'sd78823;
    data[10161] = -'sd60238;
    data[10162] =  'sd69857;
    data[10163] = -'sd2524;
    data[10164] = -'sd17668;
    data[10165] =  'sd40165;
    data[10166] = -'sd46527;
    data[10167] =  'sd1993;
    data[10168] =  'sd13951;
    data[10169] = -'sd66184;
    data[10170] =  'sd28235;
    data[10171] =  'sd33804;
    data[10172] =  'sd72787;
    data[10173] =  'sd17986;
    data[10174] = -'sd37939;
    data[10175] =  'sd62109;
    data[10176] = -'sd56760;
    data[10177] = -'sd69638;
    data[10178] =  'sd4057;
    data[10179] =  'sd28399;
    data[10180] =  'sd34952;
    data[10181] =  'sd80823;
    data[10182] =  'sd74238;
    data[10183] =  'sd28143;
    data[10184] =  'sd33160;
    data[10185] =  'sd68279;
    data[10186] = -'sd13570;
    data[10187] =  'sd68851;
    data[10188] = -'sd9566;
    data[10189] = -'sd66962;
    data[10190] =  'sd22789;
    data[10191] = -'sd4318;
    data[10192] = -'sd30226;
    data[10193] = -'sd47741;
    data[10194] = -'sd6505;
    data[10195] = -'sd45535;
    data[10196] =  'sd8937;
    data[10197] =  'sd62559;
    data[10198] = -'sd53610;
    data[10199] = -'sd47588;
    data[10200] = -'sd5434;
    data[10201] = -'sd38038;
    data[10202] =  'sd61416;
    data[10203] = -'sd61611;
    data[10204] =  'sd60246;
    data[10205] = -'sd69801;
    data[10206] =  'sd2916;
    data[10207] =  'sd20412;
    data[10208] = -'sd20957;
    data[10209] =  'sd17142;
    data[10210] = -'sd43847;
    data[10211] =  'sd20753;
    data[10212] = -'sd18570;
    data[10213] =  'sd33851;
    data[10214] =  'sd73116;
    data[10215] =  'sd20289;
    data[10216] = -'sd21818;
    data[10217] =  'sd11115;
    data[10218] =  'sd77805;
    data[10219] =  'sd53112;
    data[10220] =  'sd44102;
    data[10221] = -'sd18968;
    data[10222] =  'sd31065;
    data[10223] =  'sd53614;
    data[10224] =  'sd47616;
    data[10225] =  'sd5630;
    data[10226] =  'sd39410;
    data[10227] = -'sd51812;
    data[10228] = -'sd35002;
    data[10229] = -'sd81173;
    data[10230] = -'sd76688;
    data[10231] = -'sd45293;
    data[10232] =  'sd10631;
    data[10233] =  'sd74417;
    data[10234] =  'sd29396;
    data[10235] =  'sd41931;
    data[10236] = -'sd34165;
    data[10237] = -'sd75314;
    data[10238] = -'sd35675;
    data[10239] =  'sd77957;
    data[10240] =  'sd54176;
    data[10241] =  'sd51550;
    data[10242] =  'sd33168;
    data[10243] =  'sd68335;
    data[10244] = -'sd13178;
    data[10245] =  'sd71595;
    data[10246] =  'sd9642;
    data[10247] =  'sd67494;
    data[10248] = -'sd19065;
    data[10249] =  'sd30386;
    data[10250] =  'sd48861;
    data[10251] =  'sd14345;
    data[10252] = -'sd63426;
    data[10253] =  'sd47541;
    data[10254] =  'sd5105;
    data[10255] =  'sd35735;
    data[10256] = -'sd77537;
    data[10257] = -'sd51236;
    data[10258] = -'sd30970;
    data[10259] = -'sd52949;
    data[10260] = -'sd42961;
    data[10261] =  'sd26955;
    data[10262] =  'sd24844;
    data[10263] =  'sd10067;
    data[10264] =  'sd70469;
    data[10265] =  'sd1760;
    data[10266] =  'sd12320;
    data[10267] = -'sd77601;
    data[10268] = -'sd51684;
    data[10269] = -'sd34106;
    data[10270] = -'sd74901;
    data[10271] = -'sd32784;
    data[10272] = -'sd65647;
    data[10273] =  'sd31994;
    data[10274] =  'sd60117;
    data[10275] = -'sd70704;
    data[10276] = -'sd3405;
    data[10277] = -'sd23835;
    data[10278] = -'sd3004;
    data[10279] = -'sd21028;
    data[10280] =  'sd16645;
    data[10281] = -'sd47326;
    data[10282] = -'sd3600;
    data[10283] = -'sd25200;
    data[10284] = -'sd12559;
    data[10285] =  'sd75928;
    data[10286] =  'sd39973;
    data[10287] = -'sd47871;
    data[10288] = -'sd7415;
    data[10289] = -'sd51905;
    data[10290] = -'sd35653;
    data[10291] =  'sd78111;
    data[10292] =  'sd55254;
    data[10293] =  'sd59096;
    data[10294] = -'sd77851;
    data[10295] = -'sd53434;
    data[10296] = -'sd46356;
    data[10297] =  'sd3190;
    data[10298] =  'sd22330;
    data[10299] = -'sd7531;
    data[10300] = -'sd52717;
    data[10301] = -'sd41337;
    data[10302] =  'sd38323;
    data[10303] = -'sd59421;
    data[10304] =  'sd75576;
    data[10305] =  'sd37509;
    data[10306] = -'sd65119;
    data[10307] =  'sd35690;
    data[10308] = -'sd77852;
    data[10309] = -'sd53441;
    data[10310] = -'sd46405;
    data[10311] =  'sd2847;
    data[10312] =  'sd19929;
    data[10313] = -'sd24338;
    data[10314] = -'sd6525;
    data[10315] = -'sd45675;
    data[10316] =  'sd7957;
    data[10317] =  'sd55699;
    data[10318] =  'sd62211;
    data[10319] = -'sd56046;
    data[10320] = -'sd64640;
    data[10321] =  'sd39043;
    data[10322] = -'sd54381;
    data[10323] = -'sd52985;
    data[10324] = -'sd43213;
    data[10325] =  'sd25191;
    data[10326] =  'sd12496;
    data[10327] = -'sd76369;
    data[10328] = -'sd43060;
    data[10329] =  'sd26262;
    data[10330] =  'sd19993;
    data[10331] = -'sd23890;
    data[10332] = -'sd3389;
    data[10333] = -'sd23723;
    data[10334] = -'sd2220;
    data[10335] = -'sd15540;
    data[10336] =  'sd55061;
    data[10337] =  'sd57745;
    data[10338] =  'sd76533;
    data[10339] =  'sd44208;
    data[10340] = -'sd18226;
    data[10341] =  'sd36259;
    data[10342] = -'sd73869;
    data[10343] = -'sd25560;
    data[10344] = -'sd15079;
    data[10345] =  'sd58288;
    data[10346] =  'sd80334;
    data[10347] =  'sd70815;
    data[10348] =  'sd4182;
    data[10349] =  'sd29274;
    data[10350] =  'sd41077;
    data[10351] = -'sd40143;
    data[10352] =  'sd46681;
    data[10353] = -'sd915;
    data[10354] = -'sd6405;
    data[10355] = -'sd44835;
    data[10356] =  'sd13837;
    data[10357] = -'sd66982;
    data[10358] =  'sd22649;
    data[10359] = -'sd5298;
    data[10360] = -'sd37086;
    data[10361] =  'sd68080;
    data[10362] = -'sd14963;
    data[10363] =  'sd59100;
    data[10364] = -'sd77823;
    data[10365] = -'sd53238;
    data[10366] = -'sd44984;
    data[10367] =  'sd12794;
    data[10368] = -'sd74283;
    data[10369] = -'sd28458;
    data[10370] = -'sd35365;
    data[10371] =  'sd80127;
    data[10372] =  'sd69366;
    data[10373] = -'sd5961;
    data[10374] = -'sd41727;
    data[10375] =  'sd35593;
    data[10376] = -'sd78531;
    data[10377] = -'sd58194;
    data[10378] = -'sd79676;
    data[10379] = -'sd66209;
    data[10380] =  'sd28060;
    data[10381] =  'sd32579;
    data[10382] =  'sd64212;
    data[10383] = -'sd42039;
    data[10384] =  'sd33409;
    data[10385] =  'sd70022;
    data[10386] = -'sd1369;
    data[10387] = -'sd9583;
    data[10388] = -'sd67081;
    data[10389] =  'sd21956;
    data[10390] = -'sd10149;
    data[10391] = -'sd71043;
    data[10392] = -'sd5778;
    data[10393] = -'sd40446;
    data[10394] =  'sd44560;
    data[10395] = -'sd15762;
    data[10396] =  'sd53507;
    data[10397] =  'sd46867;
    data[10398] =  'sd387;
    data[10399] =  'sd2709;
    data[10400] =  'sd18963;
    data[10401] = -'sd31100;
    data[10402] = -'sd53859;
    data[10403] = -'sd49331;
    data[10404] = -'sd17635;
    data[10405] =  'sd40396;
    data[10406] = -'sd44910;
    data[10407] =  'sd13312;
    data[10408] = -'sd70657;
    data[10409] = -'sd3076;
    data[10410] = -'sd21532;
    data[10411] =  'sd13117;
    data[10412] = -'sd72022;
    data[10413] = -'sd12631;
    data[10414] =  'sd75424;
    data[10415] =  'sd36445;
    data[10416] = -'sd72567;
    data[10417] = -'sd16446;
    data[10418] =  'sd48719;
    data[10419] =  'sd13351;
    data[10420] = -'sd70384;
    data[10421] = -'sd1165;
    data[10422] = -'sd8155;
    data[10423] = -'sd57085;
    data[10424] = -'sd71913;
    data[10425] = -'sd11868;
    data[10426] =  'sd80765;
    data[10427] =  'sd73832;
    data[10428] =  'sd25301;
    data[10429] =  'sd13266;
    data[10430] = -'sd70979;
    data[10431] = -'sd5330;
    data[10432] = -'sd37310;
    data[10433] =  'sd66512;
    data[10434] = -'sd25939;
    data[10435] = -'sd17732;
    data[10436] =  'sd39717;
    data[10437] = -'sd49663;
    data[10438] = -'sd19959;
    data[10439] =  'sd24128;
    data[10440] =  'sd5055;
    data[10441] =  'sd35385;
    data[10442] = -'sd79987;
    data[10443] = -'sd68386;
    data[10444] =  'sd12821;
    data[10445] = -'sd74094;
    data[10446] = -'sd27135;
    data[10447] = -'sd26104;
    data[10448] = -'sd18887;
    data[10449] =  'sd31632;
    data[10450] =  'sd57583;
    data[10451] =  'sd75399;
    data[10452] =  'sd36270;
    data[10453] = -'sd73792;
    data[10454] = -'sd25021;
    data[10455] = -'sd11306;
    data[10456] = -'sd79142;
    data[10457] = -'sd62471;
    data[10458] =  'sd54226;
    data[10459] =  'sd51900;
    data[10460] =  'sd35618;
    data[10461] = -'sd78356;
    data[10462] = -'sd56969;
    data[10463] = -'sd71101;
    data[10464] = -'sd6184;
    data[10465] = -'sd43288;
    data[10466] =  'sd24666;
    data[10467] =  'sd8821;
    data[10468] =  'sd61747;
    data[10469] = -'sd59294;
    data[10470] =  'sd76465;
    data[10471] =  'sd43732;
    data[10472] = -'sd21558;
    data[10473] =  'sd12935;
    data[10474] = -'sd73296;
    data[10475] = -'sd21549;
    data[10476] =  'sd12998;
    data[10477] = -'sd72855;
    data[10478] = -'sd18462;
    data[10479] =  'sd34607;
    data[10480] =  'sd78408;
    data[10481] =  'sd57333;
    data[10482] =  'sd73649;
    data[10483] =  'sd24020;
    data[10484] =  'sd4299;
    data[10485] =  'sd30093;
    data[10486] =  'sd46810;
    data[10487] = -'sd12;
    data[10488] = -'sd84;
    data[10489] = -'sd588;
    data[10490] = -'sd4116;
    data[10491] = -'sd28812;
    data[10492] = -'sd37843;
    data[10493] =  'sd62781;
    data[10494] = -'sd52056;
    data[10495] = -'sd36710;
    data[10496] =  'sd70712;
    data[10497] =  'sd3461;
    data[10498] =  'sd24227;
    data[10499] =  'sd5748;
    data[10500] =  'sd40236;
    data[10501] = -'sd46030;
    data[10502] =  'sd5472;
    data[10503] =  'sd38304;
    data[10504] = -'sd59554;
    data[10505] =  'sd74645;
    data[10506] =  'sd30992;
    data[10507] =  'sd53103;
    data[10508] =  'sd44039;
    data[10509] = -'sd19409;
    data[10510] =  'sd27978;
    data[10511] =  'sd32005;
    data[10512] =  'sd60194;
    data[10513] = -'sd70165;
    data[10514] =  'sd368;
    data[10515] =  'sd2576;
    data[10516] =  'sd18032;
    data[10517] = -'sd37617;
    data[10518] =  'sd64363;
    data[10519] = -'sd40982;
    data[10520] =  'sd40808;
    data[10521] = -'sd42026;
    data[10522] =  'sd33500;
    data[10523] =  'sd70659;
    data[10524] =  'sd3090;
    data[10525] =  'sd21630;
    data[10526] = -'sd12431;
    data[10527] =  'sd76824;
    data[10528] =  'sd46245;
    data[10529] = -'sd3967;
    data[10530] = -'sd27769;
    data[10531] = -'sd30542;
    data[10532] = -'sd49953;
    data[10533] = -'sd21989;
    data[10534] =  'sd9918;
    data[10535] =  'sd69426;
    data[10536] = -'sd5541;
    data[10537] = -'sd38787;
    data[10538] =  'sd56173;
    data[10539] =  'sd65529;
    data[10540] = -'sd32820;
    data[10541] = -'sd65899;
    data[10542] =  'sd30230;
    data[10543] =  'sd47769;
    data[10544] =  'sd6701;
    data[10545] =  'sd46907;
    data[10546] =  'sd667;
    data[10547] =  'sd4669;
    data[10548] =  'sd32683;
    data[10549] =  'sd64940;
    data[10550] = -'sd36943;
    data[10551] =  'sd69081;
    data[10552] = -'sd7956;
    data[10553] = -'sd55692;
    data[10554] = -'sd62162;
    data[10555] =  'sd56389;
    data[10556] =  'sd67041;
    data[10557] = -'sd22236;
    data[10558] =  'sd8189;
    data[10559] =  'sd57323;
    data[10560] =  'sd73579;
    data[10561] =  'sd23530;
    data[10562] =  'sd869;
    data[10563] =  'sd6083;
    data[10564] =  'sd42581;
    data[10565] = -'sd29615;
    data[10566] = -'sd43464;
    data[10567] =  'sd23434;
    data[10568] =  'sd197;
    data[10569] =  'sd1379;
    data[10570] =  'sd9653;
    data[10571] =  'sd67571;
    data[10572] = -'sd18526;
    data[10573] =  'sd34159;
    data[10574] =  'sd75272;
    data[10575] =  'sd35381;
    data[10576] = -'sd80015;
    data[10577] = -'sd68582;
    data[10578] =  'sd11449;
    data[10579] =  'sd80143;
    data[10580] =  'sd69478;
    data[10581] = -'sd5177;
    data[10582] = -'sd36239;
    data[10583] =  'sd74009;
    data[10584] =  'sd26540;
    data[10585] =  'sd21939;
    data[10586] = -'sd10268;
    data[10587] = -'sd71876;
    data[10588] = -'sd11609;
    data[10589] = -'sd81263;
    data[10590] = -'sd77318;
    data[10591] = -'sd49703;
    data[10592] = -'sd20239;
    data[10593] =  'sd22168;
    data[10594] = -'sd8665;
    data[10595] = -'sd60655;
    data[10596] =  'sd66938;
    data[10597] = -'sd22957;
    data[10598] =  'sd3142;
    data[10599] =  'sd21994;
    data[10600] = -'sd9883;
    data[10601] = -'sd69181;
    data[10602] =  'sd7256;
    data[10603] =  'sd50792;
    data[10604] =  'sd27862;
    data[10605] =  'sd31193;
    data[10606] =  'sd54510;
    data[10607] =  'sd53888;
    data[10608] =  'sd49534;
    data[10609] =  'sd19056;
    data[10610] = -'sd30449;
    data[10611] = -'sd49302;
    data[10612] = -'sd17432;
    data[10613] =  'sd41817;
    data[10614] = -'sd34963;
    data[10615] = -'sd80900;
    data[10616] = -'sd74777;
    data[10617] = -'sd31916;
    data[10618] = -'sd59571;
    data[10619] =  'sd74526;
    data[10620] =  'sd30159;
    data[10621] =  'sd47272;
    data[10622] =  'sd3222;
    data[10623] =  'sd22554;
    data[10624] = -'sd5963;
    data[10625] = -'sd41741;
    data[10626] =  'sd35495;
    data[10627] = -'sd79217;
    data[10628] = -'sd62996;
    data[10629] =  'sd50551;
    data[10630] =  'sd26175;
    data[10631] =  'sd19384;
    data[10632] = -'sd28153;
    data[10633] = -'sd33230;
    data[10634] = -'sd68769;
    data[10635] =  'sd10140;
    data[10636] =  'sd70980;
    data[10637] =  'sd5337;
    data[10638] =  'sd37359;
    data[10639] = -'sd66169;
    data[10640] =  'sd28340;
    data[10641] =  'sd34539;
    data[10642] =  'sd77932;
    data[10643] =  'sd54001;
    data[10644] =  'sd50325;
    data[10645] =  'sd24593;
    data[10646] =  'sd8310;
    data[10647] =  'sd58170;
    data[10648] =  'sd79508;
    data[10649] =  'sd65033;
    data[10650] = -'sd36292;
    data[10651] =  'sd73638;
    data[10652] =  'sd23943;
    data[10653] =  'sd3760;
    data[10654] =  'sd26320;
    data[10655] =  'sd20399;
    data[10656] = -'sd21048;
    data[10657] =  'sd16505;
    data[10658] = -'sd48306;
    data[10659] = -'sd10460;
    data[10660] = -'sd73220;
    data[10661] = -'sd21017;
    data[10662] =  'sd16722;
    data[10663] = -'sd46787;
    data[10664] =  'sd173;
    data[10665] =  'sd1211;
    data[10666] =  'sd8477;
    data[10667] =  'sd59339;
    data[10668] = -'sd76150;
    data[10669] = -'sd41527;
    data[10670] =  'sd36993;
    data[10671] = -'sd68731;
    data[10672] =  'sd10406;
    data[10673] =  'sd72842;
    data[10674] =  'sd18371;
    data[10675] = -'sd35244;
    data[10676] =  'sd80974;
    data[10677] =  'sd75295;
    data[10678] =  'sd35542;
    data[10679] = -'sd78888;
    data[10680] = -'sd60693;
    data[10681] =  'sd66672;
    data[10682] = -'sd24819;
    data[10683] = -'sd9892;
    data[10684] = -'sd69244;
    data[10685] =  'sd6815;
    data[10686] =  'sd47705;
    data[10687] =  'sd6253;
    data[10688] =  'sd43771;
    data[10689] = -'sd21285;
    data[10690] =  'sd14846;
    data[10691] = -'sd59919;
    data[10692] =  'sd72090;
    data[10693] =  'sd13107;
    data[10694] = -'sd72092;
    data[10695] = -'sd13121;
    data[10696] =  'sd71994;
    data[10697] =  'sd12435;
    data[10698] = -'sd76796;
    data[10699] = -'sd46049;
    data[10700] =  'sd5339;
    data[10701] =  'sd37373;
    data[10702] = -'sd66071;
    data[10703] =  'sd29026;
    data[10704] =  'sd39341;
    data[10705] = -'sd52295;
    data[10706] = -'sd38383;
    data[10707] =  'sd59001;
    data[10708] = -'sd78516;
    data[10709] = -'sd58089;
    data[10710] = -'sd78941;
    data[10711] = -'sd61064;
    data[10712] =  'sd64075;
    data[10713] = -'sd42998;
    data[10714] =  'sd26696;
    data[10715] =  'sd23031;
    data[10716] = -'sd2624;
    data[10717] = -'sd18368;
    data[10718] =  'sd35265;
    data[10719] = -'sd80827;
    data[10720] = -'sd74266;
    data[10721] = -'sd28339;
    data[10722] = -'sd34532;
    data[10723] = -'sd77883;
    data[10724] = -'sd53658;
    data[10725] = -'sd47924;
    data[10726] = -'sd7786;
    data[10727] = -'sd54502;
    data[10728] = -'sd53832;
    data[10729] = -'sd49142;
    data[10730] = -'sd16312;
    data[10731] =  'sd49657;
    data[10732] =  'sd19917;
    data[10733] = -'sd24422;
    data[10734] = -'sd7113;
    data[10735] = -'sd49791;
    data[10736] = -'sd20855;
    data[10737] =  'sd17856;
    data[10738] = -'sd38849;
    data[10739] =  'sd55739;
    data[10740] =  'sd62491;
    data[10741] = -'sd54086;
    data[10742] = -'sd50920;
    data[10743] = -'sd28758;
    data[10744] = -'sd37465;
    data[10745] =  'sd65427;
    data[10746] = -'sd33534;
    data[10747] = -'sd70897;
    data[10748] = -'sd4756;
    data[10749] = -'sd33292;
    data[10750] = -'sd69203;
    data[10751] =  'sd7102;
    data[10752] =  'sd49714;
    data[10753] =  'sd20316;
    data[10754] = -'sd21629;
    data[10755] =  'sd12438;
    data[10756] = -'sd76775;
    data[10757] = -'sd45902;
    data[10758] =  'sd6368;
    data[10759] =  'sd44576;
    data[10760] = -'sd15650;
    data[10761] =  'sd54291;
    data[10762] =  'sd52355;
    data[10763] =  'sd38803;
    data[10764] = -'sd56061;
    data[10765] = -'sd64745;
    data[10766] =  'sd38308;
    data[10767] = -'sd59526;
    data[10768] =  'sd74841;
    data[10769] =  'sd32364;
    data[10770] =  'sd62707;
    data[10771] = -'sd52574;
    data[10772] = -'sd40336;
    data[10773] =  'sd45330;
    data[10774] = -'sd10372;
    data[10775] = -'sd72604;
    data[10776] = -'sd16705;
    data[10777] =  'sd46906;
    data[10778] =  'sd660;
    data[10779] =  'sd4620;
    data[10780] =  'sd32340;
    data[10781] =  'sd62539;
    data[10782] = -'sd53750;
    data[10783] = -'sd48568;
    data[10784] = -'sd12294;
    data[10785] =  'sd77783;
    data[10786] =  'sd52958;
    data[10787] =  'sd43024;
    data[10788] = -'sd26514;
    data[10789] = -'sd21757;
    data[10790] =  'sd11542;
    data[10791] =  'sd80794;
    data[10792] =  'sd74035;
    data[10793] =  'sd26722;
    data[10794] =  'sd23213;
    data[10795] = -'sd1350;
    data[10796] = -'sd9450;
    data[10797] = -'sd66150;
    data[10798] =  'sd28473;
    data[10799] =  'sd35470;
    data[10800] = -'sd79392;
    data[10801] = -'sd64221;
    data[10802] =  'sd41976;
    data[10803] = -'sd33850;
    data[10804] = -'sd73109;
    data[10805] = -'sd20240;
    data[10806] =  'sd22161;
    data[10807] = -'sd8714;
    data[10808] = -'sd60998;
    data[10809] =  'sd64537;
    data[10810] = -'sd39764;
    data[10811] =  'sd49334;
    data[10812] =  'sd17656;
    data[10813] = -'sd40249;
    data[10814] =  'sd45939;
    data[10815] = -'sd6109;
    data[10816] = -'sd42763;
    data[10817] =  'sd28341;
    data[10818] =  'sd34546;
    data[10819] =  'sd77981;
    data[10820] =  'sd54344;
    data[10821] =  'sd52726;
    data[10822] =  'sd41400;
    data[10823] = -'sd37882;
    data[10824] =  'sd62508;
    data[10825] = -'sd53967;
    data[10826] = -'sd50087;
    data[10827] = -'sd22927;
    data[10828] =  'sd3352;
    data[10829] =  'sd23464;
    data[10830] =  'sd407;
    data[10831] =  'sd2849;
    data[10832] =  'sd19943;
    data[10833] = -'sd24240;
    data[10834] = -'sd5839;
    data[10835] = -'sd40873;
    data[10836] =  'sd41571;
    data[10837] = -'sd36685;
    data[10838] =  'sd70887;
    data[10839] =  'sd4686;
    data[10840] =  'sd32802;
    data[10841] =  'sd65773;
    data[10842] = -'sd31112;
    data[10843] = -'sd53943;
    data[10844] = -'sd49919;
    data[10845] = -'sd21751;
    data[10846] =  'sd11584;
    data[10847] =  'sd81088;
    data[10848] =  'sd76093;
    data[10849] =  'sd41128;
    data[10850] = -'sd39786;
    data[10851] =  'sd49180;
    data[10852] =  'sd16578;
    data[10853] = -'sd47795;
    data[10854] = -'sd6883;
    data[10855] = -'sd48181;
    data[10856] = -'sd9585;
    data[10857] = -'sd67095;
    data[10858] =  'sd21858;
    data[10859] = -'sd10835;
    data[10860] = -'sd75845;
    data[10861] = -'sd39392;
    data[10862] =  'sd51938;
    data[10863] =  'sd35884;
    data[10864] = -'sd76494;
    data[10865] = -'sd43935;
    data[10866] =  'sd20137;
    data[10867] = -'sd22882;
    data[10868] =  'sd3667;
    data[10869] =  'sd25669;
    data[10870] =  'sd15842;
    data[10871] = -'sd52947;
    data[10872] = -'sd42947;
    data[10873] =  'sd27053;
    data[10874] =  'sd25530;
    data[10875] =  'sd14869;
    data[10876] = -'sd59758;
    data[10877] =  'sd73217;
    data[10878] =  'sd20996;
    data[10879] = -'sd16869;
    data[10880] =  'sd45758;
    data[10881] = -'sd7376;
    data[10882] = -'sd51632;
    data[10883] = -'sd33742;
    data[10884] = -'sd72353;
    data[10885] = -'sd14948;
    data[10886] =  'sd59205;
    data[10887] = -'sd77088;
    data[10888] = -'sd48093;
    data[10889] = -'sd8969;
    data[10890] = -'sd62783;
    data[10891] =  'sd52042;
    data[10892] =  'sd36612;
    data[10893] = -'sd71398;
    data[10894] = -'sd8263;
    data[10895] = -'sd57841;
    data[10896] = -'sd77205;
    data[10897] = -'sd48912;
    data[10898] = -'sd14702;
    data[10899] =  'sd60927;
    data[10900] = -'sd65034;
    data[10901] =  'sd36285;
    data[10902] = -'sd73687;
    data[10903] = -'sd24286;
    data[10904] = -'sd6161;
    data[10905] = -'sd43127;
    data[10906] =  'sd25793;
    data[10907] =  'sd16710;
    data[10908] = -'sd46871;
    data[10909] = -'sd415;
    data[10910] = -'sd2905;
    data[10911] = -'sd20335;
    data[10912] =  'sd21496;
    data[10913] = -'sd13369;
    data[10914] =  'sd70258;
    data[10915] =  'sd283;
    data[10916] =  'sd1981;
    data[10917] =  'sd13867;
    data[10918] = -'sd66772;
    data[10919] =  'sd24119;
    data[10920] =  'sd4992;
    data[10921] =  'sd34944;
    data[10922] =  'sd80767;
    data[10923] =  'sd73846;
    data[10924] =  'sd25399;
    data[10925] =  'sd13952;
    data[10926] = -'sd66177;
    data[10927] =  'sd28284;
    data[10928] =  'sd34147;
    data[10929] =  'sd75188;
    data[10930] =  'sd34793;
    data[10931] =  'sd79710;
    data[10932] =  'sd66447;
    data[10933] = -'sd26394;
    data[10934] = -'sd20917;
    data[10935] =  'sd17422;
    data[10936] = -'sd41887;
    data[10937] =  'sd34473;
    data[10938] =  'sd77470;
    data[10939] =  'sd50767;
    data[10940] =  'sd27687;
    data[10941] =  'sd29968;
    data[10942] =  'sd45935;
    data[10943] = -'sd6137;
    data[10944] = -'sd42959;
    data[10945] =  'sd26969;
    data[10946] =  'sd24942;
    data[10947] =  'sd10753;
    data[10948] =  'sd75271;
    data[10949] =  'sd35374;
    data[10950] = -'sd80064;
    data[10951] = -'sd68925;
    data[10952] =  'sd9048;
    data[10953] =  'sd63336;
    data[10954] = -'sd48171;
    data[10955] = -'sd9515;
    data[10956] = -'sd66605;
    data[10957] =  'sd25288;
    data[10958] =  'sd13175;
    data[10959] = -'sd71616;
    data[10960] = -'sd9789;
    data[10961] = -'sd68523;
    data[10962] =  'sd11862;
    data[10963] = -'sd80807;
    data[10964] = -'sd74126;
    data[10965] = -'sd27359;
    data[10966] = -'sd27672;
    data[10967] = -'sd29863;
    data[10968] = -'sd45200;
    data[10969] =  'sd11282;
    data[10970] =  'sd78974;
    data[10971] =  'sd61295;
    data[10972] = -'sd62458;
    data[10973] =  'sd54317;
    data[10974] =  'sd52537;
    data[10975] =  'sd40077;
    data[10976] = -'sd47143;
    data[10977] = -'sd2319;
    data[10978] = -'sd16233;
    data[10979] =  'sd50210;
    data[10980] =  'sd23788;
    data[10981] =  'sd2675;
    data[10982] =  'sd18725;
    data[10983] = -'sd32766;
    data[10984] = -'sd65521;
    data[10985] =  'sd32876;
    data[10986] =  'sd66291;
    data[10987] = -'sd27486;
    data[10988] = -'sd28561;
    data[10989] = -'sd36086;
    data[10990] =  'sd75080;
    data[10991] =  'sd34037;
    data[10992] =  'sd74418;
    data[10993] =  'sd29403;
    data[10994] =  'sd41980;
    data[10995] = -'sd33822;
    data[10996] = -'sd72913;
    data[10997] = -'sd18868;
    data[10998] =  'sd31765;
    data[10999] =  'sd58514;
    data[11000] =  'sd81916;
    data[11001] =  'sd81889;
    data[11002] =  'sd81700;
    data[11003] =  'sd80377;
    data[11004] =  'sd71116;
    data[11005] =  'sd6289;
    data[11006] =  'sd44023;
    data[11007] = -'sd19521;
    data[11008] =  'sd27194;
    data[11009] =  'sd26517;
    data[11010] =  'sd21778;
    data[11011] = -'sd11395;
    data[11012] = -'sd79765;
    data[11013] = -'sd66832;
    data[11014] =  'sd23699;
    data[11015] =  'sd2052;
    data[11016] =  'sd14364;
    data[11017] = -'sd63293;
    data[11018] =  'sd48472;
    data[11019] =  'sd11622;
    data[11020] =  'sd81354;
    data[11021] =  'sd77955;
    data[11022] =  'sd54162;
    data[11023] =  'sd51452;
    data[11024] =  'sd32482;
    data[11025] =  'sd63533;
    data[11026] = -'sd46792;
    data[11027] =  'sd138;
    data[11028] =  'sd966;
    data[11029] =  'sd6762;
    data[11030] =  'sd47334;
    data[11031] =  'sd3656;
    data[11032] =  'sd25592;
    data[11033] =  'sd15303;
    data[11034] = -'sd56720;
    data[11035] = -'sd69358;
    data[11036] =  'sd6017;
    data[11037] =  'sd42119;
    data[11038] = -'sd32849;
    data[11039] = -'sd66102;
    data[11040] =  'sd28809;
    data[11041] =  'sd37822;
    data[11042] = -'sd62928;
    data[11043] =  'sd51027;
    data[11044] =  'sd29507;
    data[11045] =  'sd42708;
    data[11046] = -'sd28726;
    data[11047] = -'sd37241;
    data[11048] =  'sd66995;
    data[11049] = -'sd22558;
    data[11050] =  'sd5935;
    data[11051] =  'sd41545;
    data[11052] = -'sd36867;
    data[11053] =  'sd69613;
    data[11054] = -'sd4232;
    data[11055] = -'sd29624;
    data[11056] = -'sd43527;
    data[11057] =  'sd22993;
    data[11058] = -'sd2890;
    data[11059] = -'sd20230;
    data[11060] =  'sd22231;
    data[11061] = -'sd8224;
    data[11062] = -'sd57568;
    data[11063] = -'sd75294;
    data[11064] = -'sd35535;
    data[11065] =  'sd78937;
    data[11066] =  'sd61036;
    data[11067] = -'sd64271;
    data[11068] =  'sd41626;
    data[11069] = -'sd36300;
    data[11070] =  'sd73582;
    data[11071] =  'sd23551;
    data[11072] =  'sd1016;
    data[11073] =  'sd7112;
    data[11074] =  'sd49784;
    data[11075] =  'sd20806;
    data[11076] = -'sd18199;
    data[11077] =  'sd36448;
    data[11078] = -'sd72546;
    data[11079] = -'sd16299;
    data[11080] =  'sd49748;
    data[11081] =  'sd20554;
    data[11082] = -'sd19963;
    data[11083] =  'sd24100;
    data[11084] =  'sd4859;
    data[11085] =  'sd34013;
    data[11086] =  'sd74250;
    data[11087] =  'sd28227;
    data[11088] =  'sd33748;
    data[11089] =  'sd72395;
    data[11090] =  'sd15242;
    data[11091] = -'sd57147;
    data[11092] = -'sd72347;
    data[11093] = -'sd14906;
    data[11094] =  'sd59499;
    data[11095] = -'sd75030;
    data[11096] = -'sd33687;
    data[11097] = -'sd71968;
    data[11098] = -'sd12253;
    data[11099] =  'sd78070;
    data[11100] =  'sd54967;
    data[11101] =  'sd57087;
    data[11102] =  'sd71927;
    data[11103] =  'sd11966;
    data[11104] = -'sd80079;
    data[11105] = -'sd69030;
    data[11106] =  'sd8313;
    data[11107] =  'sd58191;
    data[11108] =  'sd79655;
    data[11109] =  'sd66062;
    data[11110] = -'sd29089;
    data[11111] = -'sd39782;
    data[11112] =  'sd49208;
    data[11113] =  'sd16774;
    data[11114] = -'sd46423;
    data[11115] =  'sd2721;
    data[11116] =  'sd19047;
    data[11117] = -'sd30512;
    data[11118] = -'sd49743;
    data[11119] = -'sd20519;
    data[11120] =  'sd20208;
    data[11121] = -'sd22385;
    data[11122] =  'sd7146;
    data[11123] =  'sd50022;
    data[11124] =  'sd22472;
    data[11125] = -'sd6537;
    data[11126] = -'sd45759;
    data[11127] =  'sd7369;
    data[11128] =  'sd51583;
    data[11129] =  'sd33399;
    data[11130] =  'sd69952;
    data[11131] = -'sd1859;
    data[11132] = -'sd13013;
    data[11133] =  'sd72750;
    data[11134] =  'sd17727;
    data[11135] = -'sd39752;
    data[11136] =  'sd49418;
    data[11137] =  'sd18244;
    data[11138] = -'sd36133;
    data[11139] =  'sd74751;
    data[11140] =  'sd31734;
    data[11141] =  'sd58297;
    data[11142] =  'sd80397;
    data[11143] =  'sd71256;
    data[11144] =  'sd7269;
    data[11145] =  'sd50883;
    data[11146] =  'sd28499;
    data[11147] =  'sd35652;
    data[11148] = -'sd78118;
    data[11149] = -'sd55303;
    data[11150] = -'sd59439;
    data[11151] =  'sd75450;
    data[11152] =  'sd36627;
    data[11153] = -'sd71293;
    data[11154] = -'sd7528;
    data[11155] = -'sd52696;
    data[11156] = -'sd41190;
    data[11157] =  'sd39352;
    data[11158] = -'sd52218;
    data[11159] = -'sd37844;
    data[11160] =  'sd62774;
    data[11161] = -'sd52105;
    data[11162] = -'sd37053;
    data[11163] =  'sd68311;
    data[11164] = -'sd13346;
    data[11165] =  'sd70419;
    data[11166] =  'sd1410;
    data[11167] =  'sd9870;
    data[11168] =  'sd69090;
    data[11169] = -'sd7893;
    data[11170] = -'sd55251;
    data[11171] = -'sd59075;
    data[11172] =  'sd77998;
    data[11173] =  'sd54463;
    data[11174] =  'sd53559;
    data[11175] =  'sd47231;
    data[11176] =  'sd2935;
    data[11177] =  'sd20545;
    data[11178] = -'sd20026;
    data[11179] =  'sd23659;
    data[11180] =  'sd1772;
    data[11181] =  'sd12404;
    data[11182] = -'sd77013;
    data[11183] = -'sd47568;
    data[11184] = -'sd5294;
    data[11185] = -'sd37058;
    data[11186] =  'sd68276;
    data[11187] = -'sd13591;
    data[11188] =  'sd68704;
    data[11189] = -'sd10595;
    data[11190] = -'sd74165;
    data[11191] = -'sd27632;
    data[11192] = -'sd29583;
    data[11193] = -'sd43240;
    data[11194] =  'sd25002;
    data[11195] =  'sd11173;
    data[11196] =  'sd78211;
    data[11197] =  'sd55954;
    data[11198] =  'sd63996;
    data[11199] = -'sd43551;
    data[11200] =  'sd22825;
    data[11201] = -'sd4066;
    data[11202] = -'sd28462;
    data[11203] = -'sd35393;
    data[11204] =  'sd79931;
    data[11205] =  'sd67994;
    data[11206] = -'sd15565;
    data[11207] =  'sd54886;
    data[11208] =  'sd56520;
    data[11209] =  'sd67958;
    data[11210] = -'sd15817;
    data[11211] =  'sd53122;
    data[11212] =  'sd44172;
    data[11213] = -'sd18478;
    data[11214] =  'sd34495;
    data[11215] =  'sd77624;
    data[11216] =  'sd51845;
    data[11217] =  'sd35233;
    data[11218] = -'sd81051;
    data[11219] = -'sd75834;
    data[11220] = -'sd39315;
    data[11221] =  'sd52477;
    data[11222] =  'sd39657;
    data[11223] = -'sd50083;
    data[11224] = -'sd22899;
    data[11225] =  'sd3548;
    data[11226] =  'sd24836;
    data[11227] =  'sd10011;
    data[11228] =  'sd70077;
    data[11229] = -'sd984;
    data[11230] = -'sd6888;
    data[11231] = -'sd48216;
    data[11232] = -'sd9830;
    data[11233] = -'sd68810;
    data[11234] =  'sd9853;
    data[11235] =  'sd68971;
    data[11236] = -'sd8726;
    data[11237] = -'sd61082;
    data[11238] =  'sd63949;
    data[11239] = -'sd43880;
    data[11240] =  'sd20522;
    data[11241] = -'sd20187;
    data[11242] =  'sd22532;
    data[11243] = -'sd6117;
    data[11244] = -'sd42819;
    data[11245] =  'sd27949;
    data[11246] =  'sd31802;
    data[11247] =  'sd58773;
    data[11248] = -'sd80112;
    data[11249] = -'sd69261;
    data[11250] =  'sd6696;
    data[11251] =  'sd46872;
    data[11252] =  'sd422;
    data[11253] =  'sd2954;
    data[11254] =  'sd20678;
    data[11255] = -'sd19095;
    data[11256] =  'sd30176;
    data[11257] =  'sd47391;
    data[11258] =  'sd4055;
    data[11259] =  'sd28385;
    data[11260] =  'sd34854;
    data[11261] =  'sd80137;
    data[11262] =  'sd69436;
    data[11263] = -'sd5471;
    data[11264] = -'sd38297;
    data[11265] =  'sd59603;
    data[11266] = -'sd74302;
    data[11267] = -'sd28591;
    data[11268] = -'sd36296;
    data[11269] =  'sd73610;
    data[11270] =  'sd23747;
    data[11271] =  'sd2388;
    data[11272] =  'sd16716;
    data[11273] = -'sd46829;
    data[11274] = -'sd121;
    data[11275] = -'sd847;
    data[11276] = -'sd5929;
    data[11277] = -'sd41503;
    data[11278] =  'sd37161;
    data[11279] = -'sd67555;
    data[11280] =  'sd18638;
    data[11281] = -'sd33375;
    data[11282] = -'sd69784;
    data[11283] =  'sd3035;
    data[11284] =  'sd21245;
    data[11285] = -'sd15126;
    data[11286] =  'sd57959;
    data[11287] =  'sd78031;
    data[11288] =  'sd54694;
    data[11289] =  'sd55176;
    data[11290] =  'sd58550;
    data[11291] = -'sd81673;
    data[11292] = -'sd80188;
    data[11293] = -'sd69793;
    data[11294] =  'sd2972;
    data[11295] =  'sd20804;
    data[11296] = -'sd18213;
    data[11297] =  'sd36350;
    data[11298] = -'sd73232;
    data[11299] = -'sd21101;
    data[11300] =  'sd16134;
    data[11301] = -'sd50903;
    data[11302] = -'sd28639;
    data[11303] = -'sd36632;
    data[11304] =  'sd71258;
    data[11305] =  'sd7283;
    data[11306] =  'sd50981;
    data[11307] =  'sd29185;
    data[11308] =  'sd40454;
    data[11309] = -'sd44504;
    data[11310] =  'sd16154;
    data[11311] = -'sd50763;
    data[11312] = -'sd27659;
    data[11313] = -'sd29772;
    data[11314] = -'sd44563;
    data[11315] =  'sd15741;
    data[11316] = -'sd53654;
    data[11317] = -'sd47896;
    data[11318] = -'sd7590;
    data[11319] = -'sd53130;
    data[11320] = -'sd44228;
    data[11321] =  'sd18086;
    data[11322] = -'sd37239;
    data[11323] =  'sd67009;
    data[11324] = -'sd22460;
    data[11325] =  'sd6621;
    data[11326] =  'sd46347;
    data[11327] = -'sd3253;
    data[11328] = -'sd22771;
    data[11329] =  'sd4444;
    data[11330] =  'sd31108;
    data[11331] =  'sd53915;
    data[11332] =  'sd49723;
    data[11333] =  'sd20379;
    data[11334] = -'sd21188;
    data[11335] =  'sd15525;
    data[11336] = -'sd55166;
    data[11337] = -'sd58480;
    data[11338] = -'sd81678;
    data[11339] = -'sd80223;
    data[11340] = -'sd70038;
    data[11341] =  'sd1257;
    data[11342] =  'sd8799;
    data[11343] =  'sd61593;
    data[11344] = -'sd60372;
    data[11345] =  'sd68919;
    data[11346] = -'sd9090;
    data[11347] = -'sd63630;
    data[11348] =  'sd46113;
    data[11349] = -'sd4891;
    data[11350] = -'sd34237;
    data[11351] = -'sd75818;
    data[11352] = -'sd39203;
    data[11353] =  'sd53261;
    data[11354] =  'sd45145;
    data[11355] = -'sd11667;
    data[11356] = -'sd81669;
    data[11357] = -'sd80160;
    data[11358] = -'sd69597;
    data[11359] =  'sd4344;
    data[11360] =  'sd30408;
    data[11361] =  'sd49015;
    data[11362] =  'sd15423;
    data[11363] = -'sd55880;
    data[11364] = -'sd63478;
    data[11365] =  'sd47177;
    data[11366] =  'sd2557;
    data[11367] =  'sd17899;
    data[11368] = -'sd38548;
    data[11369] =  'sd57846;
    data[11370] =  'sd77240;
    data[11371] =  'sd49157;
    data[11372] =  'sd16417;
    data[11373] = -'sd48922;
    data[11374] = -'sd14772;
    data[11375] =  'sd60437;
    data[11376] = -'sd68464;
    data[11377] =  'sd12275;
    data[11378] = -'sd77916;
    data[11379] = -'sd53889;
    data[11380] = -'sd49541;
    data[11381] = -'sd19105;
    data[11382] =  'sd30106;
    data[11383] =  'sd46901;
    data[11384] =  'sd625;
    data[11385] =  'sd4375;
    data[11386] =  'sd30625;
    data[11387] =  'sd50534;
    data[11388] =  'sd26056;
    data[11389] =  'sd18551;
    data[11390] = -'sd33984;
    data[11391] = -'sd74047;
    data[11392] = -'sd26806;
    data[11393] = -'sd23801;
    data[11394] = -'sd2766;
    data[11395] = -'sd19362;
    data[11396] =  'sd28307;
    data[11397] =  'sd34308;
    data[11398] =  'sd76315;
    data[11399] =  'sd42682;
    data[11400] = -'sd28908;
    data[11401] = -'sd38515;
    data[11402] =  'sd58077;
    data[11403] =  'sd78857;
    data[11404] =  'sd60476;
    data[11405] = -'sd68191;
    data[11406] =  'sd14186;
    data[11407] = -'sd64539;
    data[11408] =  'sd39750;
    data[11409] = -'sd49432;
    data[11410] = -'sd18342;
    data[11411] =  'sd35447;
    data[11412] = -'sd79553;
    data[11413] = -'sd65348;
    data[11414] =  'sd34087;
    data[11415] =  'sd74768;
    data[11416] =  'sd31853;
    data[11417] =  'sd59130;
    data[11418] = -'sd77613;
    data[11419] = -'sd51768;
    data[11420] = -'sd34694;
    data[11421] = -'sd79017;
    data[11422] = -'sd61596;
    data[11423] =  'sd60351;
    data[11424] = -'sd69066;
    data[11425] =  'sd8061;
    data[11426] =  'sd56427;
    data[11427] =  'sd67307;
    data[11428] = -'sd20374;
    data[11429] =  'sd21223;
    data[11430] = -'sd15280;
    data[11431] =  'sd56881;
    data[11432] =  'sd70485;
    data[11433] =  'sd1872;
    data[11434] =  'sd13104;
    data[11435] = -'sd72113;
    data[11436] = -'sd13268;
    data[11437] =  'sd70965;
    data[11438] =  'sd5232;
    data[11439] =  'sd36624;
    data[11440] = -'sd71314;
    data[11441] = -'sd7675;
    data[11442] = -'sd53725;
    data[11443] = -'sd48393;
    data[11444] = -'sd11069;
    data[11445] = -'sd77483;
    data[11446] = -'sd50858;
    data[11447] = -'sd28324;
    data[11448] = -'sd34427;
    data[11449] = -'sd77148;
    data[11450] = -'sd48513;
    data[11451] = -'sd11909;
    data[11452] =  'sd80478;
    data[11453] =  'sd71823;
    data[11454] =  'sd11238;
    data[11455] =  'sd78666;
    data[11456] =  'sd59139;
    data[11457] = -'sd77550;
    data[11458] = -'sd51327;
    data[11459] = -'sd31607;
    data[11460] = -'sd57408;
    data[11461] = -'sd74174;
    data[11462] = -'sd27695;
    data[11463] = -'sd30024;
    data[11464] = -'sd46327;
    data[11465] =  'sd3393;
    data[11466] =  'sd23751;
    data[11467] =  'sd2416;
    data[11468] =  'sd16912;
    data[11469] = -'sd45457;
    data[11470] =  'sd9483;
    data[11471] =  'sd66381;
    data[11472] = -'sd26856;
    data[11473] = -'sd24151;
    data[11474] = -'sd5216;
    data[11475] = -'sd36512;
    data[11476] =  'sd72098;
    data[11477] =  'sd13163;
    data[11478] = -'sd71700;
    data[11479] = -'sd10377;
    data[11480] = -'sd72639;
    data[11481] = -'sd16950;
    data[11482] =  'sd45191;
    data[11483] = -'sd11345;
    data[11484] = -'sd79415;
    data[11485] = -'sd64382;
    data[11486] =  'sd40849;
    data[11487] = -'sd41739;
    data[11488] =  'sd35509;
    data[11489] = -'sd79119;
    data[11490] = -'sd62310;
    data[11491] =  'sd55353;
    data[11492] =  'sd59789;
    data[11493] = -'sd73000;
    data[11494] = -'sd19477;
    data[11495] =  'sd27502;
    data[11496] =  'sd28673;
    data[11497] =  'sd36870;
    data[11498] = -'sd69592;
    data[11499] =  'sd4379;
    data[11500] =  'sd30653;
    data[11501] =  'sd50730;
    data[11502] =  'sd27428;
    data[11503] =  'sd28155;
    data[11504] =  'sd33244;
    data[11505] =  'sd68867;
    data[11506] = -'sd9454;
    data[11507] = -'sd66178;
    data[11508] =  'sd28277;
    data[11509] =  'sd34098;
    data[11510] =  'sd74845;
    data[11511] =  'sd32392;
    data[11512] =  'sd62903;
    data[11513] = -'sd51202;
    data[11514] = -'sd30732;
    data[11515] = -'sd51283;
    data[11516] = -'sd31299;
    data[11517] = -'sd55252;
    data[11518] = -'sd59082;
    data[11519] =  'sd77949;
    data[11520] =  'sd54120;
    data[11521] =  'sd51158;
    data[11522] =  'sd30424;
    data[11523] =  'sd49127;
    data[11524] =  'sd16207;
    data[11525] = -'sd50392;
    data[11526] = -'sd25062;
    data[11527] = -'sd11593;
    data[11528] = -'sd81151;
    data[11529] = -'sd76534;
    data[11530] = -'sd44215;
    data[11531] =  'sd18177;
    data[11532] = -'sd36602;
    data[11533] =  'sd71468;
    data[11534] =  'sd8753;
    data[11535] =  'sd61271;
    data[11536] = -'sd62626;
    data[11537] =  'sd53141;
    data[11538] =  'sd44305;
    data[11539] = -'sd17547;
    data[11540] =  'sd41012;
    data[11541] = -'sd40598;
    data[11542] =  'sd43496;
    data[11543] = -'sd23210;
    data[11544] =  'sd1371;
    data[11545] =  'sd9597;
    data[11546] =  'sd67179;
    data[11547] = -'sd21270;
    data[11548] =  'sd14951;
    data[11549] = -'sd59184;
    data[11550] =  'sd77235;
    data[11551] =  'sd49122;
    data[11552] =  'sd16172;
    data[11553] = -'sd50637;
    data[11554] = -'sd26777;
    data[11555] = -'sd23598;
    data[11556] = -'sd1345;
    data[11557] = -'sd9415;
    data[11558] = -'sd65905;
    data[11559] =  'sd30188;
    data[11560] =  'sd47475;
    data[11561] =  'sd4643;
    data[11562] =  'sd32501;
    data[11563] =  'sd63666;
    data[11564] = -'sd45861;
    data[11565] =  'sd6655;
    data[11566] =  'sd46585;
    data[11567] = -'sd1587;
    data[11568] = -'sd11109;
    data[11569] = -'sd77763;
    data[11570] = -'sd52818;
    data[11571] = -'sd42044;
    data[11572] =  'sd33374;
    data[11573] =  'sd69777;
    data[11574] = -'sd3084;
    data[11575] = -'sd21588;
    data[11576] =  'sd12725;
    data[11577] = -'sd74766;
    data[11578] = -'sd31839;
    data[11579] = -'sd59032;
    data[11580] =  'sd78299;
    data[11581] =  'sd56570;
    data[11582] =  'sd68308;
    data[11583] = -'sd13367;
    data[11584] =  'sd70272;
    data[11585] =  'sd381;
    data[11586] =  'sd2667;
    data[11587] =  'sd18669;
    data[11588] = -'sd33158;
    data[11589] = -'sd68265;
    data[11590] =  'sd13668;
    data[11591] = -'sd68165;
    data[11592] =  'sd14368;
    data[11593] = -'sd63265;
    data[11594] =  'sd48668;
    data[11595] =  'sd12994;
    data[11596] = -'sd72883;
    data[11597] = -'sd18658;
    data[11598] =  'sd33235;
    data[11599] =  'sd68804;
    data[11600] = -'sd9895;
    data[11601] = -'sd69265;
    data[11602] =  'sd6668;
    data[11603] =  'sd46676;
    data[11604] = -'sd950;
    data[11605] = -'sd6650;
    data[11606] = -'sd46550;
    data[11607] =  'sd1832;
    data[11608] =  'sd12824;
    data[11609] = -'sd74073;
    data[11610] = -'sd26988;
    data[11611] = -'sd25075;
    data[11612] = -'sd11684;
    data[11613] = -'sd81788;
    data[11614] = -'sd80993;
    data[11615] = -'sd75428;
    data[11616] = -'sd36473;
    data[11617] =  'sd72371;
    data[11618] =  'sd15074;
    data[11619] = -'sd58323;
    data[11620] = -'sd80579;
    data[11621] = -'sd72530;
    data[11622] = -'sd16187;
    data[11623] =  'sd50532;
    data[11624] =  'sd26042;
    data[11625] =  'sd18453;
    data[11626] = -'sd34670;
    data[11627] = -'sd78849;
    data[11628] = -'sd60420;
    data[11629] =  'sd68583;
    data[11630] = -'sd11442;
    data[11631] = -'sd80094;
    data[11632] = -'sd69135;
    data[11633] =  'sd7578;
    data[11634] =  'sd53046;
    data[11635] =  'sd43640;
    data[11636] = -'sd22202;
    data[11637] =  'sd8427;
    data[11638] =  'sd58989;
    data[11639] = -'sd78600;
    data[11640] = -'sd58677;
    data[11641] =  'sd80784;
    data[11642] =  'sd73965;
    data[11643] =  'sd26232;
    data[11644] =  'sd19783;
    data[11645] = -'sd25360;
    data[11646] = -'sd13679;
    data[11647] =  'sd68088;
    data[11648] = -'sd14907;
    data[11649] =  'sd59492;
    data[11650] = -'sd75079;
    data[11651] = -'sd34030;
    data[11652] = -'sd74369;
    data[11653] = -'sd29060;
    data[11654] = -'sd39579;
    data[11655] =  'sd50629;
    data[11656] =  'sd26721;
    data[11657] =  'sd23206;
    data[11658] = -'sd1399;
    data[11659] = -'sd9793;
    data[11660] = -'sd68551;
    data[11661] =  'sd11666;
    data[11662] =  'sd81662;
    data[11663] =  'sd80111;
    data[11664] =  'sd69254;
    data[11665] = -'sd6745;
    data[11666] = -'sd47215;
    data[11667] = -'sd2823;
    data[11668] = -'sd19761;
    data[11669] =  'sd25514;
    data[11670] =  'sd14757;
    data[11671] = -'sd60542;
    data[11672] =  'sd67729;
    data[11673] = -'sd17420;
    data[11674] =  'sd41901;
    data[11675] = -'sd34375;
    data[11676] = -'sd76784;
    data[11677] = -'sd45965;
    data[11678] =  'sd5927;
    data[11679] =  'sd41489;
    data[11680] = -'sd37259;
    data[11681] =  'sd66869;
    data[11682] = -'sd23440;
    data[11683] = -'sd239;
    data[11684] = -'sd1673;
    data[11685] = -'sd11711;
    data[11686] =  'sd81864;
    data[11687] =  'sd81525;
    data[11688] =  'sd79152;
    data[11689] =  'sd62541;
    data[11690] = -'sd53736;
    data[11691] = -'sd48470;
    data[11692] = -'sd11608;
    data[11693] = -'sd81256;
    data[11694] = -'sd77269;
    data[11695] = -'sd49360;
    data[11696] = -'sd17838;
    data[11697] =  'sd38975;
    data[11698] = -'sd54857;
    data[11699] = -'sd56317;
    data[11700] = -'sd66537;
    data[11701] =  'sd25764;
    data[11702] =  'sd16507;
    data[11703] = -'sd48292;
    data[11704] = -'sd10362;
    data[11705] = -'sd72534;
    data[11706] = -'sd16215;
    data[11707] =  'sd50336;
    data[11708] =  'sd24670;
    data[11709] =  'sd8849;
    data[11710] =  'sd61943;
    data[11711] = -'sd57922;
    data[11712] = -'sd77772;
    data[11713] = -'sd52881;
    data[11714] = -'sd42485;
    data[11715] =  'sd30287;
    data[11716] =  'sd48168;
    data[11717] =  'sd9494;
    data[11718] =  'sd66458;
    data[11719] = -'sd26317;
    data[11720] = -'sd20378;
    data[11721] =  'sd21195;
    data[11722] = -'sd15476;
    data[11723] =  'sd55509;
    data[11724] =  'sd60881;
    data[11725] = -'sd65356;
    data[11726] =  'sd34031;
    data[11727] =  'sd74376;
    data[11728] =  'sd29109;
    data[11729] =  'sd39922;
    data[11730] = -'sd48228;
    data[11731] = -'sd9914;
    data[11732] = -'sd69398;
    data[11733] =  'sd5737;
    data[11734] =  'sd40159;
    data[11735] = -'sd46569;
    data[11736] =  'sd1699;
    data[11737] =  'sd11893;
    data[11738] = -'sd80590;
    data[11739] = -'sd72607;
    data[11740] = -'sd16726;
    data[11741] =  'sd46759;
    data[11742] = -'sd369;
    data[11743] = -'sd2583;
    data[11744] = -'sd18081;
    data[11745] =  'sd37274;
    data[11746] = -'sd66764;
    data[11747] =  'sd24175;
    data[11748] =  'sd5384;
    data[11749] =  'sd37688;
    data[11750] = -'sd63866;
    data[11751] =  'sd44461;
    data[11752] = -'sd16455;
    data[11753] =  'sd48656;
    data[11754] =  'sd12910;
    data[11755] = -'sd73471;
    data[11756] = -'sd22774;
    data[11757] =  'sd4423;
    data[11758] =  'sd30961;
    data[11759] =  'sd52886;
    data[11760] =  'sd42520;
    data[11761] = -'sd30042;
    data[11762] = -'sd46453;
    data[11763] =  'sd2511;
    data[11764] =  'sd17577;
    data[11765] = -'sd40802;
    data[11766] =  'sd42068;
    data[11767] = -'sd33206;
    data[11768] = -'sd68601;
    data[11769] =  'sd11316;
    data[11770] =  'sd79212;
    data[11771] =  'sd62961;
    data[11772] = -'sd50796;
    data[11773] = -'sd27890;
    data[11774] = -'sd31389;
    data[11775] = -'sd55882;
    data[11776] = -'sd63492;
    data[11777] =  'sd47079;
    data[11778] =  'sd1871;
    data[11779] =  'sd13097;
    data[11780] = -'sd72162;
    data[11781] = -'sd13611;
    data[11782] =  'sd68564;
    data[11783] = -'sd11575;
    data[11784] = -'sd81025;
    data[11785] = -'sd75652;
    data[11786] = -'sd38041;
    data[11787] =  'sd61395;
    data[11788] = -'sd61758;
    data[11789] =  'sd59217;
    data[11790] = -'sd77004;
    data[11791] = -'sd47505;
    data[11792] = -'sd4853;
    data[11793] = -'sd33971;
    data[11794] = -'sd73956;
    data[11795] = -'sd26169;
    data[11796] = -'sd19342;
    data[11797] =  'sd28447;
    data[11798] =  'sd35288;
    data[11799] = -'sd80666;
    data[11800] = -'sd73139;
    data[11801] = -'sd20450;
    data[11802] =  'sd20691;
    data[11803] = -'sd19004;
    data[11804] =  'sd30813;
    data[11805] =  'sd51850;
    data[11806] =  'sd35268;
    data[11807] = -'sd80806;
    data[11808] = -'sd74119;
    data[11809] = -'sd27310;
    data[11810] = -'sd27329;
    data[11811] = -'sd27462;
    data[11812] = -'sd28393;
    data[11813] = -'sd34910;
    data[11814] = -'sd80529;
    data[11815] = -'sd72180;
    data[11816] = -'sd13737;
    data[11817] =  'sd67682;
    data[11818] = -'sd17749;
    data[11819] =  'sd39598;
    data[11820] = -'sd50496;
    data[11821] = -'sd25790;
    data[11822] = -'sd16689;
    data[11823] =  'sd47018;
    data[11824] =  'sd1444;
    data[11825] =  'sd10108;
    data[11826] =  'sd70756;
    data[11827] =  'sd3769;
    data[11828] =  'sd26383;
    data[11829] =  'sd20840;
    data[11830] = -'sd17961;
    data[11831] =  'sd38114;
    data[11832] = -'sd60884;
    data[11833] =  'sd65335;
    data[11834] = -'sd34178;
    data[11835] = -'sd75405;
    data[11836] = -'sd36312;
    data[11837] =  'sd73498;
    data[11838] =  'sd22963;
    data[11839] = -'sd3100;
    data[11840] = -'sd21700;
    data[11841] =  'sd11941;
    data[11842] = -'sd80254;
    data[11843] = -'sd70255;
    data[11844] = -'sd262;
    data[11845] = -'sd1834;
    data[11846] = -'sd12838;
    data[11847] =  'sd73975;
    data[11848] =  'sd26302;
    data[11849] =  'sd20273;
    data[11850] = -'sd21930;
    data[11851] =  'sd10331;
    data[11852] =  'sd72317;
    data[11853] =  'sd14696;
    data[11854] = -'sd60969;
    data[11855] =  'sd64740;
    data[11856] = -'sd38343;
    data[11857] =  'sd59281;
    data[11858] = -'sd76556;
    data[11859] = -'sd44369;
    data[11860] =  'sd17099;
    data[11861] = -'sd44148;
    data[11862] =  'sd18646;
    data[11863] = -'sd33319;
    data[11864] = -'sd69392;
    data[11865] =  'sd5779;
    data[11866] =  'sd40453;
    data[11867] = -'sd44511;
    data[11868] =  'sd16105;
    data[11869] = -'sd51106;
    data[11870] = -'sd30060;
    data[11871] = -'sd46579;
    data[11872] =  'sd1629;
    data[11873] =  'sd11403;
    data[11874] =  'sd79821;
    data[11875] =  'sd67224;
    data[11876] = -'sd20955;
    data[11877] =  'sd17156;
    data[11878] = -'sd43749;
    data[11879] =  'sd21439;
    data[11880] = -'sd13768;
    data[11881] =  'sd67465;
    data[11882] = -'sd19268;
    data[11883] =  'sd28965;
    data[11884] =  'sd38914;
    data[11885] = -'sd55284;
    data[11886] = -'sd59306;
    data[11887] =  'sd76381;
    data[11888] =  'sd43144;
    data[11889] = -'sd25674;
    data[11890] = -'sd15877;
    data[11891] =  'sd52702;
    data[11892] =  'sd41232;
    data[11893] = -'sd39058;
    data[11894] =  'sd54276;
    data[11895] =  'sd52250;
    data[11896] =  'sd38068;
    data[11897] = -'sd61206;
    data[11898] =  'sd63081;
    data[11899] = -'sd49956;
    data[11900] = -'sd22010;
    data[11901] =  'sd9771;
    data[11902] =  'sd68397;
    data[11903] = -'sd12744;
    data[11904] =  'sd74633;
    data[11905] =  'sd30908;
    data[11906] =  'sd52515;
    data[11907] =  'sd39923;
    data[11908] = -'sd48221;
    data[11909] = -'sd9865;
    data[11910] = -'sd69055;
    data[11911] =  'sd8138;
    data[11912] =  'sd56966;
    data[11913] =  'sd71080;
    data[11914] =  'sd6037;
    data[11915] =  'sd42259;
    data[11916] = -'sd31869;
    data[11917] = -'sd59242;
    data[11918] =  'sd76829;
    data[11919] =  'sd46280;
    data[11920] = -'sd3722;
    data[11921] = -'sd26054;
    data[11922] = -'sd18537;
    data[11923] =  'sd34082;
    data[11924] =  'sd74733;
    data[11925] =  'sd31608;
    data[11926] =  'sd57415;
    data[11927] =  'sd74223;
    data[11928] =  'sd28038;
    data[11929] =  'sd32425;
    data[11930] =  'sd63134;
    data[11931] = -'sd49585;
    data[11932] = -'sd19413;
    data[11933] =  'sd27950;
    data[11934] =  'sd31809;
    data[11935] =  'sd58822;
    data[11936] = -'sd79769;
    data[11937] = -'sd66860;
    data[11938] =  'sd23503;
    data[11939] =  'sd680;
    data[11940] =  'sd4760;
    data[11941] =  'sd33320;
    data[11942] =  'sd69399;
    data[11943] = -'sd5730;
    data[11944] = -'sd40110;
    data[11945] =  'sd46912;
    data[11946] =  'sd702;
    data[11947] =  'sd4914;
    data[11948] =  'sd34398;
    data[11949] =  'sd76945;
    data[11950] =  'sd47092;
    data[11951] =  'sd1962;
    data[11952] =  'sd13734;
    data[11953] = -'sd67703;
    data[11954] =  'sd17602;
    data[11955] = -'sd40627;
    data[11956] =  'sd43293;
    data[11957] = -'sd24631;
    data[11958] = -'sd8576;
    data[11959] = -'sd60032;
    data[11960] =  'sd71299;
    data[11961] =  'sd7570;
    data[11962] =  'sd52990;
    data[11963] =  'sd43248;
    data[11964] = -'sd24946;
    data[11965] = -'sd10781;
    data[11966] = -'sd75467;
    data[11967] = -'sd36746;
    data[11968] =  'sd70460;
    data[11969] =  'sd1697;
    data[11970] =  'sd11879;
    data[11971] = -'sd80688;
    data[11972] = -'sd73293;
    data[11973] = -'sd21528;
    data[11974] =  'sd13145;
    data[11975] = -'sd71826;
    data[11976] = -'sd11259;
    data[11977] = -'sd78813;
    data[11978] = -'sd60168;
    data[11979] =  'sd70347;
    data[11980] =  'sd906;
    data[11981] =  'sd6342;
    data[11982] =  'sd44394;
    data[11983] = -'sd16924;
    data[11984] =  'sd45373;
    data[11985] = -'sd10071;
    data[11986] = -'sd70497;
    data[11987] = -'sd1956;
    data[11988] = -'sd13692;
    data[11989] =  'sd67997;
    data[11990] = -'sd15544;
    data[11991] =  'sd55033;
    data[11992] =  'sd57549;
    data[11993] =  'sd75161;
    data[11994] =  'sd34604;
    data[11995] =  'sd78387;
    data[11996] =  'sd57186;
    data[11997] =  'sd72620;
    data[11998] =  'sd16817;
    data[11999] = -'sd46122;
    data[12000] =  'sd4828;
    data[12001] =  'sd33796;
    data[12002] =  'sd72731;
    data[12003] =  'sd17594;
    data[12004] = -'sd40683;
    data[12005] =  'sd42901;
    data[12006] = -'sd27375;
    data[12007] = -'sd27784;
    data[12008] = -'sd30647;
    data[12009] = -'sd50688;
    data[12010] = -'sd27134;
    data[12011] = -'sd26097;
    data[12012] = -'sd18838;
    data[12013] =  'sd31975;
    data[12014] =  'sd59984;
    data[12015] = -'sd71635;
    data[12016] = -'sd9922;
    data[12017] = -'sd69454;
    data[12018] =  'sd5345;
    data[12019] =  'sd37415;
    data[12020] = -'sd65777;
    data[12021] =  'sd31084;
    data[12022] =  'sd53747;
    data[12023] =  'sd48547;
    data[12024] =  'sd12147;
    data[12025] = -'sd78812;
    data[12026] = -'sd60161;
    data[12027] =  'sd70396;
    data[12028] =  'sd1249;
    data[12029] =  'sd8743;
    data[12030] =  'sd61201;
    data[12031] = -'sd63116;
    data[12032] =  'sd49711;
    data[12033] =  'sd20295;
    data[12034] = -'sd21776;
    data[12035] =  'sd11409;
    data[12036] =  'sd79863;
    data[12037] =  'sd67518;
    data[12038] = -'sd18897;
    data[12039] =  'sd31562;
    data[12040] =  'sd57093;
    data[12041] =  'sd71969;
    data[12042] =  'sd12260;
    data[12043] = -'sd78021;
    data[12044] = -'sd54624;
    data[12045] = -'sd54686;
    data[12046] = -'sd55120;
    data[12047] = -'sd58158;
    data[12048] = -'sd79424;
    data[12049] = -'sd64445;
    data[12050] =  'sd40408;
    data[12051] = -'sd44826;
    data[12052] =  'sd13900;
    data[12053] = -'sd66541;
    data[12054] =  'sd25736;
    data[12055] =  'sd16311;
    data[12056] = -'sd49664;
    data[12057] = -'sd19966;
    data[12058] =  'sd24079;
    data[12059] =  'sd4712;
    data[12060] =  'sd32984;
    data[12061] =  'sd67047;
    data[12062] = -'sd22194;
    data[12063] =  'sd8483;
    data[12064] =  'sd59381;
    data[12065] = -'sd75856;
    data[12066] = -'sd39469;
    data[12067] =  'sd51399;
    data[12068] =  'sd32111;
    data[12069] =  'sd60936;
    data[12070] = -'sd64971;
    data[12071] =  'sd36726;
    data[12072] = -'sd70600;
    data[12073] = -'sd2677;
    data[12074] = -'sd18739;
    data[12075] =  'sd32668;
    data[12076] =  'sd64835;
    data[12077] = -'sd37678;
    data[12078] =  'sd63936;
    data[12079] = -'sd43971;
    data[12080] =  'sd19885;
    data[12081] = -'sd24646;
    data[12082] = -'sd8681;
    data[12083] = -'sd60767;
    data[12084] =  'sd66154;
    data[12085] = -'sd28445;
    data[12086] = -'sd35274;
    data[12087] =  'sd80764;
    data[12088] =  'sd73825;
    data[12089] =  'sd25252;
    data[12090] =  'sd12923;
    data[12091] = -'sd73380;
    data[12092] = -'sd22137;
    data[12093] =  'sd8882;
    data[12094] =  'sd62174;
    data[12095] = -'sd56305;
    data[12096] = -'sd66453;
    data[12097] =  'sd26352;
    data[12098] =  'sd20623;
    data[12099] = -'sd19480;
    data[12100] =  'sd27481;
    data[12101] =  'sd28526;
    data[12102] =  'sd35841;
    data[12103] = -'sd76795;
    data[12104] = -'sd46042;
    data[12105] =  'sd5388;
    data[12106] =  'sd37716;
    data[12107] = -'sd63670;
    data[12108] =  'sd45833;
    data[12109] = -'sd6851;
    data[12110] = -'sd47957;
    data[12111] = -'sd8017;
    data[12112] = -'sd56119;
    data[12113] = -'sd65151;
    data[12114] =  'sd35466;
    data[12115] = -'sd79420;
    data[12116] = -'sd64417;
    data[12117] =  'sd40604;
    data[12118] = -'sd43454;
    data[12119] =  'sd23504;
    data[12120] =  'sd687;
    data[12121] =  'sd4809;
    data[12122] =  'sd33663;
    data[12123] =  'sd71800;
    data[12124] =  'sd11077;
    data[12125] =  'sd77539;
    data[12126] =  'sd51250;
    data[12127] =  'sd31068;
    data[12128] =  'sd53635;
    data[12129] =  'sd47763;
    data[12130] =  'sd6659;
    data[12131] =  'sd46613;
    data[12132] = -'sd1391;
    data[12133] = -'sd9737;
    data[12134] = -'sd68159;
    data[12135] =  'sd14410;
    data[12136] = -'sd62971;
    data[12137] =  'sd50726;
    data[12138] =  'sd27400;
    data[12139] =  'sd27959;
    data[12140] =  'sd31872;
    data[12141] =  'sd59263;
    data[12142] = -'sd76682;
    data[12143] = -'sd45251;
    data[12144] =  'sd10925;
    data[12145] =  'sd76475;
    data[12146] =  'sd43802;
    data[12147] = -'sd21068;
    data[12148] =  'sd16365;
    data[12149] = -'sd49286;
    data[12150] = -'sd17320;
    data[12151] =  'sd42601;
    data[12152] = -'sd29475;
    data[12153] = -'sd42484;
    data[12154] =  'sd30294;
    data[12155] =  'sd48217;
    data[12156] =  'sd9837;
    data[12157] =  'sd68859;
    data[12158] = -'sd9510;
    data[12159] = -'sd66570;
    data[12160] =  'sd25533;
    data[12161] =  'sd14890;
    data[12162] = -'sd59611;
    data[12163] =  'sd74246;
    data[12164] =  'sd28199;
    data[12165] =  'sd33552;
    data[12166] =  'sd71023;
    data[12167] =  'sd5638;
    data[12168] =  'sd39466;
    data[12169] = -'sd51420;
    data[12170] = -'sd32258;
    data[12171] = -'sd61965;
    data[12172] =  'sd57768;
    data[12173] =  'sd76694;
    data[12174] =  'sd45335;
    data[12175] = -'sd10337;
    data[12176] = -'sd72359;
    data[12177] = -'sd14990;
    data[12178] =  'sd58911;
    data[12179] = -'sd79146;
    data[12180] = -'sd62499;
    data[12181] =  'sd54030;
    data[12182] =  'sd50528;
    data[12183] =  'sd26014;
    data[12184] =  'sd18257;
    data[12185] = -'sd36042;
    data[12186] =  'sd75388;
    data[12187] =  'sd36193;
    data[12188] = -'sd74331;
    data[12189] = -'sd28794;
    data[12190] = -'sd37717;
    data[12191] =  'sd63663;
    data[12192] = -'sd45882;
    data[12193] =  'sd6508;
    data[12194] =  'sd45556;
    data[12195] = -'sd8790;
    data[12196] = -'sd61530;
    data[12197] =  'sd60813;
    data[12198] = -'sd65832;
    data[12199] =  'sd30699;
    data[12200] =  'sd51052;
    data[12201] =  'sd29682;
    data[12202] =  'sd43933;
    data[12203] = -'sd20151;
    data[12204] =  'sd22784;
    data[12205] = -'sd4353;
    data[12206] = -'sd30471;
    data[12207] = -'sd49456;
    data[12208] = -'sd18510;
    data[12209] =  'sd34271;
    data[12210] =  'sd76056;
    data[12211] =  'sd40869;
    data[12212] = -'sd41599;
    data[12213] =  'sd36489;
    data[12214] = -'sd72259;
    data[12215] = -'sd14290;
    data[12216] =  'sd63811;
    data[12217] = -'sd44846;
    data[12218] =  'sd13760;
    data[12219] = -'sd67521;
    data[12220] =  'sd18876;
    data[12221] = -'sd31709;
    data[12222] = -'sd58122;
    data[12223] = -'sd79172;
    data[12224] = -'sd62681;
    data[12225] =  'sd52756;
    data[12226] =  'sd41610;
    data[12227] = -'sd36412;
    data[12228] =  'sd72798;
    data[12229] =  'sd18063;
    data[12230] = -'sd37400;
    data[12231] =  'sd65882;
    data[12232] = -'sd30349;
    data[12233] = -'sd48602;
    data[12234] = -'sd12532;
    data[12235] =  'sd76117;
    data[12236] =  'sd41296;
    data[12237] = -'sd38610;
    data[12238] =  'sd57412;
    data[12239] =  'sd74202;
    data[12240] =  'sd27891;
    data[12241] =  'sd31396;
    data[12242] =  'sd55931;
    data[12243] =  'sd63835;
    data[12244] = -'sd44678;
    data[12245] =  'sd14936;
    data[12246] = -'sd59289;
    data[12247] =  'sd76500;
    data[12248] =  'sd43977;
    data[12249] = -'sd19843;
    data[12250] =  'sd24940;
    data[12251] =  'sd10739;
    data[12252] =  'sd75173;
    data[12253] =  'sd34688;
    data[12254] =  'sd78975;
    data[12255] =  'sd61302;
    data[12256] = -'sd62409;
    data[12257] =  'sd54660;
    data[12258] =  'sd54938;
    data[12259] =  'sd56884;
    data[12260] =  'sd70506;
    data[12261] =  'sd2019;
    data[12262] =  'sd14133;
    data[12263] = -'sd64910;
    data[12264] =  'sd37153;
    data[12265] = -'sd67611;
    data[12266] =  'sd18246;
    data[12267] = -'sd36119;
    data[12268] =  'sd74849;
    data[12269] =  'sd32420;
    data[12270] =  'sd63099;
    data[12271] = -'sd49830;
    data[12272] = -'sd21128;
    data[12273] =  'sd15945;
    data[12274] = -'sd52226;
    data[12275] = -'sd37900;
    data[12276] =  'sd62382;
    data[12277] = -'sd54849;
    data[12278] = -'sd56261;
    data[12279] = -'sd66145;
    data[12280] =  'sd28508;
    data[12281] =  'sd35715;
    data[12282] = -'sd77677;
    data[12283] = -'sd52216;
    data[12284] = -'sd37830;
    data[12285] =  'sd62872;
    data[12286] = -'sd51419;
    data[12287] = -'sd32251;
    data[12288] = -'sd61916;
    data[12289] =  'sd58111;
    data[12290] =  'sd79095;
    data[12291] =  'sd62142;
    data[12292] = -'sd56529;
    data[12293] = -'sd68021;
    data[12294] =  'sd15376;
    data[12295] = -'sd56209;
    data[12296] = -'sd65781;
    data[12297] =  'sd31056;
    data[12298] =  'sd53551;
    data[12299] =  'sd47175;
    data[12300] =  'sd2543;
    data[12301] =  'sd17801;
    data[12302] = -'sd39234;
    data[12303] =  'sd53044;
    data[12304] =  'sd43626;
    data[12305] = -'sd22300;
    data[12306] =  'sd7741;
    data[12307] =  'sd54187;
    data[12308] =  'sd51627;
    data[12309] =  'sd33707;
    data[12310] =  'sd72108;
    data[12311] =  'sd13233;
    data[12312] = -'sd71210;
    data[12313] = -'sd6947;
    data[12314] = -'sd48629;
    data[12315] = -'sd12721;
    data[12316] =  'sd74794;
    data[12317] =  'sd32035;
    data[12318] =  'sd60404;
    data[12319] = -'sd68695;
    data[12320] =  'sd10658;
    data[12321] =  'sd74606;
    data[12322] =  'sd30719;
    data[12323] =  'sd51192;
    data[12324] =  'sd30662;
    data[12325] =  'sd50793;
    data[12326] =  'sd27869;
    data[12327] =  'sd31242;
    data[12328] =  'sd54853;
    data[12329] =  'sd56289;
    data[12330] =  'sd66341;
    data[12331] = -'sd27136;
    data[12332] = -'sd26111;
    data[12333] = -'sd18936;
    data[12334] =  'sd31289;
    data[12335] =  'sd55182;
    data[12336] =  'sd58592;
    data[12337] = -'sd81379;
    data[12338] = -'sd78130;
    data[12339] = -'sd55387;
    data[12340] = -'sd60027;
    data[12341] =  'sd71334;
    data[12342] =  'sd7815;
    data[12343] =  'sd54705;
    data[12344] =  'sd55253;
    data[12345] =  'sd59089;
    data[12346] = -'sd77900;
    data[12347] = -'sd53777;
    data[12348] = -'sd48757;
    data[12349] = -'sd13617;
    data[12350] =  'sd68522;
    data[12351] = -'sd11869;
    data[12352] =  'sd80758;
    data[12353] =  'sd73783;
    data[12354] =  'sd24958;
    data[12355] =  'sd10865;
    data[12356] =  'sd76055;
    data[12357] =  'sd40862;
    data[12358] = -'sd41648;
    data[12359] =  'sd36146;
    data[12360] = -'sd74660;
    data[12361] = -'sd31097;
    data[12362] = -'sd53838;
    data[12363] = -'sd49184;
    data[12364] = -'sd16606;
    data[12365] =  'sd47599;
    data[12366] =  'sd5511;
    data[12367] =  'sd38577;
    data[12368] = -'sd57643;
    data[12369] = -'sd75819;
    data[12370] = -'sd39210;
    data[12371] =  'sd53212;
    data[12372] =  'sd44802;
    data[12373] = -'sd14068;
    data[12374] =  'sd65365;
    data[12375] = -'sd33968;
    data[12376] = -'sd73935;
    data[12377] = -'sd26022;
    data[12378] = -'sd18313;
    data[12379] =  'sd35650;
    data[12380] = -'sd78132;
    data[12381] = -'sd55401;
    data[12382] = -'sd60125;
    data[12383] =  'sd70648;
    data[12384] =  'sd3013;
    data[12385] =  'sd21091;
    data[12386] = -'sd16204;
    data[12387] =  'sd50413;
    data[12388] =  'sd25209;
    data[12389] =  'sd12622;
    data[12390] = -'sd75487;
    data[12391] = -'sd36886;
    data[12392] =  'sd69480;
    data[12393] = -'sd5163;
    data[12394] = -'sd36141;
    data[12395] =  'sd74695;
    data[12396] =  'sd31342;
    data[12397] =  'sd55553;
    data[12398] =  'sd61189;
    data[12399] = -'sd63200;
    data[12400] =  'sd49123;
    data[12401] =  'sd16179;
    data[12402] = -'sd50588;
    data[12403] = -'sd26434;
    data[12404] = -'sd21197;
    data[12405] =  'sd15462;
    data[12406] = -'sd55607;
    data[12407] = -'sd61567;
    data[12408] =  'sd60554;
    data[12409] = -'sd67645;
    data[12410] =  'sd18008;
    data[12411] = -'sd37785;
    data[12412] =  'sd63187;
    data[12413] = -'sd49214;
    data[12414] = -'sd16816;
    data[12415] =  'sd46129;
    data[12416] = -'sd4779;
    data[12417] = -'sd33453;
    data[12418] = -'sd70330;
    data[12419] = -'sd787;
    data[12420] = -'sd5509;
    data[12421] = -'sd38563;
    data[12422] =  'sd57741;
    data[12423] =  'sd76505;
    data[12424] =  'sd44012;
    data[12425] = -'sd19598;
    data[12426] =  'sd26655;
    data[12427] =  'sd22744;
    data[12428] = -'sd4633;
    data[12429] = -'sd32431;
    data[12430] = -'sd63176;
    data[12431] =  'sd49291;
    data[12432] =  'sd17355;
    data[12433] = -'sd42356;
    data[12434] =  'sd31190;
    data[12435] =  'sd54489;
    data[12436] =  'sd53741;
    data[12437] =  'sd48505;
    data[12438] =  'sd11853;
    data[12439] = -'sd80870;
    data[12440] = -'sd74567;
    data[12441] = -'sd30446;
    data[12442] = -'sd49281;
    data[12443] = -'sd17285;
    data[12444] =  'sd42846;
    data[12445] = -'sd27760;
    data[12446] = -'sd30479;
    data[12447] = -'sd49512;
    data[12448] = -'sd18902;
    data[12449] =  'sd31527;
    data[12450] =  'sd56848;
    data[12451] =  'sd70254;
    data[12452] =  'sd255;
    data[12453] =  'sd1785;
    data[12454] =  'sd12495;
    data[12455] = -'sd76376;
    data[12456] = -'sd43109;
    data[12457] =  'sd25919;
    data[12458] =  'sd17592;
    data[12459] = -'sd40697;
    data[12460] =  'sd42803;
    data[12461] = -'sd28061;
    data[12462] = -'sd32586;
    data[12463] = -'sd64261;
    data[12464] =  'sd41696;
    data[12465] = -'sd35810;
    data[12466] =  'sd77012;
    data[12467] =  'sd47561;
    data[12468] =  'sd5245;
    data[12469] =  'sd36715;
    data[12470] = -'sd70677;
    data[12471] = -'sd3216;
    data[12472] = -'sd22512;
    data[12473] =  'sd6257;
    data[12474] =  'sd43799;
    data[12475] = -'sd21089;
    data[12476] =  'sd16218;
    data[12477] = -'sd50315;
    data[12478] = -'sd24523;
    data[12479] = -'sd7820;
    data[12480] = -'sd54740;
    data[12481] = -'sd55498;
    data[12482] = -'sd60804;
    data[12483] =  'sd65895;
    data[12484] = -'sd30258;
    data[12485] = -'sd47965;
    data[12486] = -'sd8073;
    data[12487] = -'sd56511;
    data[12488] = -'sd67895;
    data[12489] =  'sd16258;
    data[12490] = -'sd50035;
    data[12491] = -'sd22563;
    data[12492] =  'sd5900;
    data[12493] =  'sd41300;
    data[12494] = -'sd38582;
    data[12495] =  'sd57608;
    data[12496] =  'sd75574;
    data[12497] =  'sd37495;
    data[12498] = -'sd65217;
    data[12499] =  'sd35004;
    data[12500] =  'sd81187;
    data[12501] =  'sd76786;
    data[12502] =  'sd45979;
    data[12503] = -'sd5829;
    data[12504] = -'sd40803;
    data[12505] =  'sd42061;
    data[12506] = -'sd33255;
    data[12507] = -'sd68944;
    data[12508] =  'sd8915;
    data[12509] =  'sd62405;
    data[12510] = -'sd54688;
    data[12511] = -'sd55134;
    data[12512] = -'sd58256;
    data[12513] = -'sd80110;
    data[12514] = -'sd69247;
    data[12515] =  'sd6794;
    data[12516] =  'sd47558;
    data[12517] =  'sd5224;
    data[12518] =  'sd36568;
    data[12519] = -'sd71706;
    data[12520] = -'sd10419;
    data[12521] = -'sd72933;
    data[12522] = -'sd19008;
    data[12523] =  'sd30785;
    data[12524] =  'sd51654;
    data[12525] =  'sd33896;
    data[12526] =  'sd73431;
    data[12527] =  'sd22494;
    data[12528] = -'sd6383;
    data[12529] = -'sd44681;
    data[12530] =  'sd14915;
    data[12531] = -'sd59436;
    data[12532] =  'sd75471;
    data[12533] =  'sd36774;
    data[12534] = -'sd70264;
    data[12535] = -'sd325;
    data[12536] = -'sd2275;
    data[12537] = -'sd15925;
    data[12538] =  'sd52366;
    data[12539] =  'sd38880;
    data[12540] = -'sd55522;
    data[12541] = -'sd60972;
    data[12542] =  'sd64719;
    data[12543] = -'sd38490;
    data[12544] =  'sd58252;
    data[12545] =  'sd80082;
    data[12546] =  'sd69051;
    data[12547] = -'sd8166;
    data[12548] = -'sd57162;
    data[12549] = -'sd72452;
    data[12550] = -'sd15641;
    data[12551] =  'sd54354;
    data[12552] =  'sd52796;
    data[12553] =  'sd41890;
    data[12554] = -'sd34452;
    data[12555] = -'sd77323;
    data[12556] = -'sd49738;
    data[12557] = -'sd20484;
    data[12558] =  'sd20453;
    data[12559] = -'sd20670;
    data[12560] =  'sd19151;
    data[12561] = -'sd29784;
    data[12562] = -'sd44647;
    data[12563] =  'sd15153;
    data[12564] = -'sd57770;
    data[12565] = -'sd76708;
    data[12566] = -'sd45433;
    data[12567] =  'sd9651;
    data[12568] =  'sd67557;
    data[12569] = -'sd18624;
    data[12570] =  'sd33473;
    data[12571] =  'sd70470;
    data[12572] =  'sd1767;
    data[12573] =  'sd12369;
    data[12574] = -'sd77258;
    data[12575] = -'sd49283;
    data[12576] = -'sd17299;
    data[12577] =  'sd42748;
    data[12578] = -'sd28446;
    data[12579] = -'sd35281;
    data[12580] =  'sd80715;
    data[12581] =  'sd73482;
    data[12582] =  'sd22851;
    data[12583] = -'sd3884;
    data[12584] = -'sd27188;
    data[12585] = -'sd26475;
    data[12586] = -'sd21484;
    data[12587] =  'sd13453;
    data[12588] = -'sd69670;
    data[12589] =  'sd3833;
    data[12590] =  'sd26831;
    data[12591] =  'sd23976;
    data[12592] =  'sd3991;
    data[12593] =  'sd27937;
    data[12594] =  'sd31718;
    data[12595] =  'sd58185;
    data[12596] =  'sd79613;
    data[12597] =  'sd65768;
    data[12598] = -'sd31147;
    data[12599] = -'sd54188;
    data[12600] = -'sd51634;
    data[12601] = -'sd33756;
    data[12602] = -'sd72451;
    data[12603] = -'sd15634;
    data[12604] =  'sd54403;
    data[12605] =  'sd53139;
    data[12606] =  'sd44291;
    data[12607] = -'sd17645;
    data[12608] =  'sd40326;
    data[12609] = -'sd45400;
    data[12610] =  'sd9882;
    data[12611] =  'sd69174;
    data[12612] = -'sd7305;
    data[12613] = -'sd51135;
    data[12614] = -'sd30263;
    data[12615] = -'sd48000;
    data[12616] = -'sd8318;
    data[12617] = -'sd58226;
    data[12618] = -'sd79900;
    data[12619] = -'sd67777;
    data[12620] =  'sd17084;
    data[12621] = -'sd44253;
    data[12622] =  'sd17911;
    data[12623] = -'sd38464;
    data[12624] =  'sd58434;
    data[12625] =  'sd81356;
    data[12626] =  'sd77969;
    data[12627] =  'sd54260;
    data[12628] =  'sd52138;
    data[12629] =  'sd37284;
    data[12630] = -'sd66694;
    data[12631] =  'sd24665;
    data[12632] =  'sd8814;
    data[12633] =  'sd61698;
    data[12634] = -'sd59637;
    data[12635] =  'sd74064;
    data[12636] =  'sd26925;
    data[12637] =  'sd24634;
    data[12638] =  'sd8597;
    data[12639] =  'sd60179;
    data[12640] = -'sd70270;
    data[12641] = -'sd367;
    data[12642] = -'sd2569;
    data[12643] = -'sd17983;
    data[12644] =  'sd37960;
    data[12645] = -'sd61962;
    data[12646] =  'sd57789;
    data[12647] =  'sd76841;
    data[12648] =  'sd46364;
    data[12649] = -'sd3134;
    data[12650] = -'sd21938;
    data[12651] =  'sd10275;
    data[12652] =  'sd71925;
    data[12653] =  'sd11952;
    data[12654] = -'sd80177;
    data[12655] = -'sd69716;
    data[12656] =  'sd3511;
    data[12657] =  'sd24577;
    data[12658] =  'sd8198;
    data[12659] =  'sd57386;
    data[12660] =  'sd74020;
    data[12661] =  'sd26617;
    data[12662] =  'sd22478;
    data[12663] = -'sd6495;
    data[12664] = -'sd45465;
    data[12665] =  'sd9427;
    data[12666] =  'sd65989;
    data[12667] = -'sd29600;
    data[12668] = -'sd43359;
    data[12669] =  'sd24169;
    data[12670] =  'sd5342;
    data[12671] =  'sd37394;
    data[12672] = -'sd65924;
    data[12673] =  'sd30055;
    data[12674] =  'sd46544;
    data[12675] = -'sd1874;
    data[12676] = -'sd13118;
    data[12677] =  'sd72015;
    data[12678] =  'sd12582;
    data[12679] = -'sd75767;
    data[12680] = -'sd38846;
    data[12681] =  'sd55760;
    data[12682] =  'sd62638;
    data[12683] = -'sd53057;
    data[12684] = -'sd43717;
    data[12685] =  'sd21663;
    data[12686] = -'sd12200;
    data[12687] =  'sd78441;
    data[12688] =  'sd57564;
    data[12689] =  'sd75266;
    data[12690] =  'sd35339;
    data[12691] = -'sd80309;
    data[12692] = -'sd70640;
    data[12693] = -'sd2957;
    data[12694] = -'sd20699;
    data[12695] =  'sd18948;
    data[12696] = -'sd31205;
    data[12697] = -'sd54594;
    data[12698] = -'sd54476;
    data[12699] = -'sd53650;
    data[12700] = -'sd47868;
    data[12701] = -'sd7394;
    data[12702] = -'sd51758;
    data[12703] = -'sd34624;
    data[12704] = -'sd78527;
    data[12705] = -'sd58166;
    data[12706] = -'sd79480;
    data[12707] = -'sd64837;
    data[12708] =  'sd37664;
    data[12709] = -'sd64034;
    data[12710] =  'sd43285;
    data[12711] = -'sd24687;
    data[12712] = -'sd8968;
    data[12713] = -'sd62776;
    data[12714] =  'sd52091;
    data[12715] =  'sd36955;
    data[12716] = -'sd68997;
    data[12717] =  'sd8544;
    data[12718] =  'sd59808;
    data[12719] = -'sd72867;
    data[12720] = -'sd18546;
    data[12721] =  'sd34019;
    data[12722] =  'sd74292;
    data[12723] =  'sd28521;
    data[12724] =  'sd35806;
    data[12725] = -'sd77040;
    data[12726] = -'sd47757;
    data[12727] = -'sd6617;
    data[12728] = -'sd46319;
    data[12729] =  'sd3449;
    data[12730] =  'sd24143;
    data[12731] =  'sd5160;
    data[12732] =  'sd36120;
    data[12733] = -'sd74842;
    data[12734] = -'sd32371;
    data[12735] = -'sd62756;
    data[12736] =  'sd52231;
    data[12737] =  'sd37935;
    data[12738] = -'sd62137;
    data[12739] =  'sd56564;
    data[12740] =  'sd68266;
    data[12741] = -'sd13661;
    data[12742] =  'sd68214;
    data[12743] = -'sd14025;
    data[12744] =  'sd65666;
    data[12745] = -'sd31861;
    data[12746] = -'sd59186;
    data[12747] =  'sd77221;
    data[12748] =  'sd49024;
    data[12749] =  'sd15486;
    data[12750] = -'sd55439;
    data[12751] = -'sd60391;
    data[12752] =  'sd68786;
    data[12753] = -'sd10021;
    data[12754] = -'sd70147;
    data[12755] =  'sd494;
    data[12756] =  'sd3458;
    data[12757] =  'sd24206;
    data[12758] =  'sd5601;
    data[12759] =  'sd39207;
    data[12760] = -'sd53233;
    data[12761] = -'sd44949;
    data[12762] =  'sd13039;
    data[12763] = -'sd72568;
    data[12764] = -'sd16453;
    data[12765] =  'sd48670;
    data[12766] =  'sd13008;
    data[12767] = -'sd72785;
    data[12768] = -'sd17972;
    data[12769] =  'sd38037;
    data[12770] = -'sd61423;
    data[12771] =  'sd61562;
    data[12772] = -'sd60589;
    data[12773] =  'sd67400;
    data[12774] = -'sd19723;
    data[12775] =  'sd25780;
    data[12776] =  'sd16619;
    data[12777] = -'sd47508;
    data[12778] = -'sd4874;
    data[12779] = -'sd34118;
    data[12780] = -'sd74985;
    data[12781] = -'sd33372;
    data[12782] = -'sd69763;
    data[12783] =  'sd3182;
    data[12784] =  'sd22274;
    data[12785] = -'sd7923;
    data[12786] = -'sd55461;
    data[12787] = -'sd60545;
    data[12788] =  'sd67708;
    data[12789] = -'sd17567;
    data[12790] =  'sd40872;
    data[12791] = -'sd41578;
    data[12792] =  'sd36636;
    data[12793] = -'sd71230;
    data[12794] = -'sd7087;
    data[12795] = -'sd49609;
    data[12796] = -'sd19581;
    data[12797] =  'sd26774;
    data[12798] =  'sd23577;
    data[12799] =  'sd1198;
    data[12800] =  'sd8386;
    data[12801] =  'sd58702;
    data[12802] = -'sd80609;
    data[12803] = -'sd72740;
    data[12804] = -'sd17657;
    data[12805] =  'sd40242;
    data[12806] = -'sd45988;
    data[12807] =  'sd5766;
    data[12808] =  'sd40362;
    data[12809] = -'sd45148;
    data[12810] =  'sd11646;
    data[12811] =  'sd81522;
    data[12812] =  'sd79131;
    data[12813] =  'sd62394;
    data[12814] = -'sd54765;
    data[12815] = -'sd55673;
    data[12816] = -'sd62029;
    data[12817] =  'sd57320;
    data[12818] =  'sd73558;
    data[12819] =  'sd23383;
    data[12820] = -'sd160;
    data[12821] = -'sd1120;
    data[12822] = -'sd7840;
    data[12823] = -'sd54880;
    data[12824] = -'sd56478;
    data[12825] = -'sd67664;
    data[12826] =  'sd17875;
    data[12827] = -'sd38716;
    data[12828] =  'sd56670;
    data[12829] =  'sd69008;
    data[12830] = -'sd8467;
    data[12831] = -'sd59269;
    data[12832] =  'sd76640;
    data[12833] =  'sd44957;
    data[12834] = -'sd12983;
    data[12835] =  'sd72960;
    data[12836] =  'sd19197;
    data[12837] = -'sd29462;
    data[12838] = -'sd42393;
    data[12839] =  'sd30931;
    data[12840] =  'sd52676;
    data[12841] =  'sd41050;
    data[12842] = -'sd40332;
    data[12843] =  'sd45358;
    data[12844] = -'sd10176;
    data[12845] = -'sd71232;
    data[12846] = -'sd7101;
    data[12847] = -'sd49707;
    data[12848] = -'sd20267;
    data[12849] =  'sd21972;
    data[12850] = -'sd10037;
    data[12851] = -'sd70259;
    data[12852] = -'sd290;
    data[12853] = -'sd2030;
    data[12854] = -'sd14210;
    data[12855] =  'sd64371;
    data[12856] = -'sd40926;
    data[12857] =  'sd41200;
    data[12858] = -'sd39282;
    data[12859] =  'sd52708;
    data[12860] =  'sd41274;
    data[12861] = -'sd38764;
    data[12862] =  'sd56334;
    data[12863] =  'sd66656;
    data[12864] = -'sd24931;
    data[12865] = -'sd10676;
    data[12866] = -'sd74732;
    data[12867] = -'sd31601;
    data[12868] = -'sd57366;
    data[12869] = -'sd73880;
    data[12870] = -'sd25637;
    data[12871] = -'sd15618;
    data[12872] =  'sd54515;
    data[12873] =  'sd53923;
    data[12874] =  'sd49779;
    data[12875] =  'sd20771;
    data[12876] = -'sd18444;
    data[12877] =  'sd34733;
    data[12878] =  'sd79290;
    data[12879] =  'sd63507;
    data[12880] = -'sd46974;
    data[12881] = -'sd1136;
    data[12882] = -'sd7952;
    data[12883] = -'sd55664;
    data[12884] = -'sd61966;
    data[12885] =  'sd57761;
    data[12886] =  'sd76645;
    data[12887] =  'sd44992;
    data[12888] = -'sd12738;
    data[12889] =  'sd74675;
    data[12890] =  'sd31202;
    data[12891] =  'sd54573;
    data[12892] =  'sd54329;
    data[12893] =  'sd52621;
    data[12894] =  'sd40665;
    data[12895] = -'sd43027;
    data[12896] =  'sd26493;
    data[12897] =  'sd21610;
    data[12898] = -'sd12571;
    data[12899] =  'sd75844;
    data[12900] =  'sd39385;
    data[12901] = -'sd51987;
    data[12902] = -'sd36227;
    data[12903] =  'sd74093;
    data[12904] =  'sd27128;
    data[12905] =  'sd26055;
    data[12906] =  'sd18544;
    data[12907] = -'sd34033;
    data[12908] = -'sd74390;
    data[12909] = -'sd29207;
    data[12910] = -'sd40608;
    data[12911] =  'sd43426;
    data[12912] = -'sd23700;
    data[12913] = -'sd2059;
    data[12914] = -'sd14413;
    data[12915] =  'sd62950;
    data[12916] = -'sd50873;
    data[12917] = -'sd28429;
    data[12918] = -'sd35162;
    data[12919] =  'sd81548;
    data[12920] =  'sd79313;
    data[12921] =  'sd63668;
    data[12922] = -'sd45847;
    data[12923] =  'sd6753;
    data[12924] =  'sd47271;
    data[12925] =  'sd3215;
    data[12926] =  'sd22505;
    data[12927] = -'sd6306;
    data[12928] = -'sd44142;
    data[12929] =  'sd18688;
    data[12930] = -'sd33025;
    data[12931] = -'sd67334;
    data[12932] =  'sd20185;
    data[12933] = -'sd22546;
    data[12934] =  'sd6019;
    data[12935] =  'sd42133;
    data[12936] = -'sd32751;
    data[12937] = -'sd65416;
    data[12938] =  'sd33611;
    data[12939] =  'sd71436;
    data[12940] =  'sd8529;
    data[12941] =  'sd59703;
    data[12942] = -'sd73602;
    data[12943] = -'sd23691;
    data[12944] = -'sd1996;
    data[12945] = -'sd13972;
    data[12946] =  'sd66037;
    data[12947] = -'sd29264;
    data[12948] = -'sd41007;
    data[12949] =  'sd40633;
    data[12950] = -'sd43251;
    data[12951] =  'sd24925;
    data[12952] =  'sd10634;
    data[12953] =  'sd74438;
    data[12954] =  'sd29543;
    data[12955] =  'sd42960;
    data[12956] = -'sd26962;
    data[12957] = -'sd24893;
    data[12958] = -'sd10410;
    data[12959] = -'sd72870;
    data[12960] = -'sd18567;
    data[12961] =  'sd33872;
    data[12962] =  'sd73263;
    data[12963] =  'sd21318;
    data[12964] = -'sd14615;
    data[12965] =  'sd61536;
    data[12966] = -'sd60771;
    data[12967] =  'sd66126;
    data[12968] = -'sd28641;
    data[12969] = -'sd36646;
    data[12970] =  'sd71160;
    data[12971] =  'sd6597;
    data[12972] =  'sd46179;
    data[12973] = -'sd4429;
    data[12974] = -'sd31003;
    data[12975] = -'sd53180;
    data[12976] = -'sd44578;
    data[12977] =  'sd15636;
    data[12978] = -'sd54389;
    data[12979] = -'sd53041;
    data[12980] = -'sd43605;
    data[12981] =  'sd22447;
    data[12982] = -'sd6712;
    data[12983] = -'sd46984;
    data[12984] = -'sd1206;
    data[12985] = -'sd8442;
    data[12986] = -'sd59094;
    data[12987] =  'sd77865;
    data[12988] =  'sd53532;
    data[12989] =  'sd47042;
    data[12990] =  'sd1612;
    data[12991] =  'sd11284;
    data[12992] =  'sd78988;
    data[12993] =  'sd61393;
    data[12994] = -'sd61772;
    data[12995] =  'sd59119;
    data[12996] = -'sd77690;
    data[12997] = -'sd52307;
    data[12998] = -'sd38467;
    data[12999] =  'sd58413;
    data[13000] =  'sd81209;
    data[13001] =  'sd76940;
    data[13002] =  'sd47057;
    data[13003] =  'sd1717;
    data[13004] =  'sd12019;
    data[13005] = -'sd79708;
    data[13006] = -'sd66433;
    data[13007] =  'sd26492;
    data[13008] =  'sd21603;
    data[13009] = -'sd12620;
    data[13010] =  'sd75501;
    data[13011] =  'sd36984;
    data[13012] = -'sd68794;
    data[13013] =  'sd9965;
    data[13014] =  'sd69755;
    data[13015] = -'sd3238;
    data[13016] = -'sd22666;
    data[13017] =  'sd5179;
    data[13018] =  'sd36253;
    data[13019] = -'sd73911;
    data[13020] = -'sd25854;
    data[13021] = -'sd17137;
    data[13022] =  'sd43882;
    data[13023] = -'sd20508;
    data[13024] =  'sd20285;
    data[13025] = -'sd21846;
    data[13026] =  'sd10919;
    data[13027] =  'sd76433;
    data[13028] =  'sd43508;
    data[13029] = -'sd23126;
    data[13030] =  'sd1959;
    data[13031] =  'sd13713;
    data[13032] = -'sd67850;
    data[13033] =  'sd16573;
    data[13034] = -'sd47830;
    data[13035] = -'sd7128;
    data[13036] = -'sd49896;
    data[13037] = -'sd21590;
    data[13038] =  'sd12711;
    data[13039] = -'sd74864;
    data[13040] = -'sd32525;
    data[13041] = -'sd63834;
    data[13042] =  'sd44685;
    data[13043] = -'sd14887;
    data[13044] =  'sd59632;
    data[13045] = -'sd74099;
    data[13046] = -'sd27170;
    data[13047] = -'sd26349;
    data[13048] = -'sd20602;
    data[13049] =  'sd19627;
    data[13050] = -'sd26452;
    data[13051] = -'sd21323;
    data[13052] =  'sd14580;
    data[13053] = -'sd61781;
    data[13054] =  'sd59056;
    data[13055] = -'sd78131;
    data[13056] = -'sd55394;
    data[13057] = -'sd60076;
    data[13058] =  'sd70991;
    data[13059] =  'sd5414;
    data[13060] =  'sd37898;
    data[13061] = -'sd62396;
    data[13062] =  'sd54751;
    data[13063] =  'sd55575;
    data[13064] =  'sd61343;
    data[13065] = -'sd62122;
    data[13066] =  'sd56669;
    data[13067] =  'sd69001;
    data[13068] = -'sd8516;
    data[13069] = -'sd59612;
    data[13070] =  'sd74239;
    data[13071] =  'sd28150;
    data[13072] =  'sd33209;
    data[13073] =  'sd68622;
    data[13074] = -'sd11169;
    data[13075] = -'sd78183;
    data[13076] = -'sd55758;
    data[13077] = -'sd62624;
    data[13078] =  'sd53155;
    data[13079] =  'sd44403;
    data[13080] = -'sd16861;
    data[13081] =  'sd45814;
    data[13082] = -'sd6984;
    data[13083] = -'sd48888;
    data[13084] = -'sd14534;
    data[13085] =  'sd62103;
    data[13086] = -'sd56802;
    data[13087] = -'sd69932;
    data[13088] =  'sd1999;
    data[13089] =  'sd13993;
    data[13090] = -'sd65890;
    data[13091] =  'sd30293;
    data[13092] =  'sd48210;
    data[13093] =  'sd9788;
    data[13094] =  'sd68516;
    data[13095] = -'sd11911;
    data[13096] =  'sd80464;
    data[13097] =  'sd71725;
    data[13098] =  'sd10552;
    data[13099] =  'sd73864;
    data[13100] =  'sd25525;
    data[13101] =  'sd14834;
    data[13102] = -'sd60003;
    data[13103] =  'sd71502;
    data[13104] =  'sd8991;
    data[13105] =  'sd62937;
    data[13106] = -'sd50964;
    data[13107] = -'sd29066;
    data[13108] = -'sd39621;
    data[13109] =  'sd50335;
    data[13110] =  'sd24663;
    data[13111] =  'sd8800;
    data[13112] =  'sd61600;
    data[13113] = -'sd60323;
    data[13114] =  'sd69262;
    data[13115] = -'sd6689;
    data[13116] = -'sd46823;
    data[13117] = -'sd79;
    data[13118] = -'sd553;
    data[13119] = -'sd3871;
    data[13120] = -'sd27097;
    data[13121] = -'sd25838;
    data[13122] = -'sd17025;
    data[13123] =  'sd44666;
    data[13124] = -'sd15020;
    data[13125] =  'sd58701;
    data[13126] = -'sd80616;
    data[13127] = -'sd72789;
    data[13128] = -'sd18000;
    data[13129] =  'sd37841;
    data[13130] = -'sd62795;
    data[13131] =  'sd51958;
    data[13132] =  'sd36024;
    data[13133] = -'sd75514;
    data[13134] = -'sd37075;
    data[13135] =  'sd68157;
    data[13136] = -'sd14424;
    data[13137] =  'sd62873;
    data[13138] = -'sd51412;
    data[13139] = -'sd32202;
    data[13140] = -'sd61573;
    data[13141] =  'sd60512;
    data[13142] = -'sd67939;
    data[13143] =  'sd15950;
    data[13144] = -'sd52191;
    data[13145] = -'sd37655;
    data[13146] =  'sd64097;
    data[13147] = -'sd42844;
    data[13148] =  'sd27774;
    data[13149] =  'sd30577;
    data[13150] =  'sd50198;
    data[13151] =  'sd23704;
    data[13152] =  'sd2087;
    data[13153] =  'sd14609;
    data[13154] = -'sd61578;
    data[13155] =  'sd60477;
    data[13156] = -'sd68184;
    data[13157] =  'sd14235;
    data[13158] = -'sd64196;
    data[13159] =  'sd42151;
    data[13160] = -'sd32625;
    data[13161] = -'sd64534;
    data[13162] =  'sd39785;
    data[13163] = -'sd49187;
    data[13164] = -'sd16627;
    data[13165] =  'sd47452;
    data[13166] =  'sd4482;
    data[13167] =  'sd31374;
    data[13168] =  'sd55777;
    data[13169] =  'sd62757;
    data[13170] = -'sd52224;
    data[13171] = -'sd37886;
    data[13172] =  'sd62480;
    data[13173] = -'sd54163;
    data[13174] = -'sd51459;
    data[13175] = -'sd32531;
    data[13176] = -'sd63876;
    data[13177] =  'sd44391;
    data[13178] = -'sd16945;
    data[13179] =  'sd45226;
    data[13180] = -'sd11100;
    data[13181] = -'sd77700;
    data[13182] = -'sd52377;
    data[13183] = -'sd38957;
    data[13184] =  'sd54983;
    data[13185] =  'sd57199;
    data[13186] =  'sd72711;
    data[13187] =  'sd17454;
    data[13188] = -'sd41663;
    data[13189] =  'sd36041;
    data[13190] = -'sd75395;
    data[13191] = -'sd36242;
    data[13192] =  'sd73988;
    data[13193] =  'sd26393;
    data[13194] =  'sd20910;
    data[13195] = -'sd17471;
    data[13196] =  'sd41544;
    data[13197] = -'sd36874;
    data[13198] =  'sd69564;
    data[13199] = -'sd4575;
    data[13200] = -'sd32025;
    data[13201] = -'sd60334;
    data[13202] =  'sd69185;
    data[13203] = -'sd7228;
    data[13204] = -'sd50596;
    data[13205] = -'sd26490;
    data[13206] = -'sd21589;
    data[13207] =  'sd12718;
    data[13208] = -'sd74815;
    data[13209] = -'sd32182;
    data[13210] = -'sd61433;
    data[13211] =  'sd61492;
    data[13212] = -'sd61079;
    data[13213] =  'sd63970;
    data[13214] = -'sd43733;
    data[13215] =  'sd21551;
    data[13216] = -'sd12984;
    data[13217] =  'sd72953;
    data[13218] =  'sd19148;
    data[13219] = -'sd29805;
    data[13220] = -'sd44794;
    data[13221] =  'sd14124;
    data[13222] = -'sd64973;
    data[13223] =  'sd36712;
    data[13224] = -'sd70698;
    data[13225] = -'sd3363;
    data[13226] = -'sd23541;
    data[13227] = -'sd946;
    data[13228] = -'sd6622;
    data[13229] = -'sd46354;
    data[13230] =  'sd3204;
    data[13231] =  'sd22428;
    data[13232] = -'sd6845;
    data[13233] = -'sd47915;
    data[13234] = -'sd7723;
    data[13235] = -'sd54061;
    data[13236] = -'sd50745;
    data[13237] = -'sd27533;
    data[13238] = -'sd28890;
    data[13239] = -'sd38389;
    data[13240] =  'sd58959;
    data[13241] = -'sd78810;
    data[13242] = -'sd60147;
    data[13243] =  'sd70494;
    data[13244] =  'sd1935;
    data[13245] =  'sd13545;
    data[13246] = -'sd69026;
    data[13247] =  'sd8341;
    data[13248] =  'sd58387;
    data[13249] =  'sd81027;
    data[13250] =  'sd75666;
    data[13251] =  'sd38139;
    data[13252] = -'sd60709;
    data[13253] =  'sd66560;
    data[13254] = -'sd25603;
    data[13255] = -'sd15380;
    data[13256] =  'sd56181;
    data[13257] =  'sd65585;
    data[13258] = -'sd32428;
    data[13259] = -'sd63155;
    data[13260] =  'sd49438;
    data[13261] =  'sd18384;
    data[13262] = -'sd35153;
    data[13263] =  'sd81611;
    data[13264] =  'sd79754;
    data[13265] =  'sd66755;
    data[13266] = -'sd24238;
    data[13267] = -'sd5825;
    data[13268] = -'sd40775;
    data[13269] =  'sd42257;
    data[13270] = -'sd31883;
    data[13271] = -'sd59340;
    data[13272] =  'sd76143;
    data[13273] =  'sd41478;
    data[13274] = -'sd37336;
    data[13275] =  'sd66330;
    data[13276] = -'sd27213;
    data[13277] = -'sd26650;
    data[13278] = -'sd22709;
    data[13279] =  'sd4878;
    data[13280] =  'sd34146;
    data[13281] =  'sd75181;
    data[13282] =  'sd34744;
    data[13283] =  'sd79367;
    data[13284] =  'sd64046;
    data[13285] = -'sd43201;
    data[13286] =  'sd25275;
    data[13287] =  'sd13084;
    data[13288] = -'sd72253;
    data[13289] = -'sd14248;
    data[13290] =  'sd64105;
    data[13291] = -'sd42788;
    data[13292] =  'sd28166;
    data[13293] =  'sd33321;
    data[13294] =  'sd69406;
    data[13295] = -'sd5681;
    data[13296] = -'sd39767;
    data[13297] =  'sd49313;
    data[13298] =  'sd17509;
    data[13299] = -'sd41278;
    data[13300] =  'sd38736;
    data[13301] = -'sd56530;
    data[13302] = -'sd68028;
    data[13303] =  'sd15327;
    data[13304] = -'sd56552;
    data[13305] = -'sd68182;
    data[13306] =  'sd14249;
    data[13307] = -'sd64098;
    data[13308] =  'sd42837;
    data[13309] = -'sd27823;
    data[13310] = -'sd30920;
    data[13311] = -'sd52599;
    data[13312] = -'sd40511;
    data[13313] =  'sd44105;
    data[13314] = -'sd18947;
    data[13315] =  'sd31212;
    data[13316] =  'sd54643;
    data[13317] =  'sd54819;
    data[13318] =  'sd56051;
    data[13319] =  'sd64675;
    data[13320] = -'sd38798;
    data[13321] =  'sd56096;
    data[13322] =  'sd64990;
    data[13323] = -'sd36593;
    data[13324] =  'sd71531;
    data[13325] =  'sd9194;
    data[13326] =  'sd64358;
    data[13327] = -'sd41017;
    data[13328] =  'sd40563;
    data[13329] = -'sd43741;
    data[13330] =  'sd21495;
    data[13331] = -'sd13376;
    data[13332] =  'sd70209;
    data[13333] = -'sd60;
    data[13334] = -'sd420;
    data[13335] = -'sd2940;
    data[13336] = -'sd20580;
    data[13337] =  'sd19781;
    data[13338] = -'sd25374;
    data[13339] = -'sd13777;
    data[13340] =  'sd67402;
    data[13341] = -'sd19709;
    data[13342] =  'sd25878;
    data[13343] =  'sd17305;
    data[13344] = -'sd42706;
    data[13345] =  'sd28740;
    data[13346] =  'sd37339;
    data[13347] = -'sd66309;
    data[13348] =  'sd27360;
    data[13349] =  'sd27679;
    data[13350] =  'sd29912;
    data[13351] =  'sd45543;
    data[13352] = -'sd8881;
    data[13353] = -'sd62167;
    data[13354] =  'sd56354;
    data[13355] =  'sd66796;
    data[13356] = -'sd23951;
    data[13357] = -'sd3816;
    data[13358] = -'sd26712;
    data[13359] = -'sd23143;
    data[13360] =  'sd1840;
    data[13361] =  'sd12880;
    data[13362] = -'sd73681;
    data[13363] = -'sd24244;
    data[13364] = -'sd5867;
    data[13365] = -'sd41069;
    data[13366] =  'sd40199;
    data[13367] = -'sd46289;
    data[13368] =  'sd3659;
    data[13369] =  'sd25613;
    data[13370] =  'sd15450;
    data[13371] = -'sd55691;
    data[13372] = -'sd62155;
    data[13373] =  'sd56438;
    data[13374] =  'sd67384;
    data[13375] = -'sd19835;
    data[13376] =  'sd24996;
    data[13377] =  'sd11131;
    data[13378] =  'sd77917;
    data[13379] =  'sd53896;
    data[13380] =  'sd49590;
    data[13381] =  'sd19448;
    data[13382] = -'sd27705;
    data[13383] = -'sd30094;
    data[13384] = -'sd46817;
    data[13385] = -'sd37;
    data[13386] = -'sd259;
    data[13387] = -'sd1813;
    data[13388] = -'sd12691;
    data[13389] =  'sd75004;
    data[13390] =  'sd33505;
    data[13391] =  'sd70694;
    data[13392] =  'sd3335;
    data[13393] =  'sd23345;
    data[13394] = -'sd426;
    data[13395] = -'sd2982;
    data[13396] = -'sd20874;
    data[13397] =  'sd17723;
    data[13398] = -'sd39780;
    data[13399] =  'sd49222;
    data[13400] =  'sd16872;
    data[13401] = -'sd45737;
    data[13402] =  'sd7523;
    data[13403] =  'sd52661;
    data[13404] =  'sd40945;
    data[13405] = -'sd41067;
    data[13406] =  'sd40213;
    data[13407] = -'sd46191;
    data[13408] =  'sd4345;
    data[13409] =  'sd30415;
    data[13410] =  'sd49064;
    data[13411] =  'sd15766;
    data[13412] = -'sd53479;
    data[13413] = -'sd46671;
    data[13414] =  'sd985;
    data[13415] =  'sd6895;
    data[13416] =  'sd48265;
    data[13417] =  'sd10173;
    data[13418] =  'sd71211;
    data[13419] =  'sd6954;
    data[13420] =  'sd48678;
    data[13421] =  'sd13064;
    data[13422] = -'sd72393;
    data[13423] = -'sd15228;
    data[13424] =  'sd57245;
    data[13425] =  'sd73033;
    data[13426] =  'sd19708;
    data[13427] = -'sd25885;
    data[13428] = -'sd17354;
    data[13429] =  'sd42363;
    data[13430] = -'sd31141;
    data[13431] = -'sd54146;
    data[13432] = -'sd51340;
    data[13433] = -'sd31698;
    data[13434] = -'sd58045;
    data[13435] = -'sd78633;
    data[13436] = -'sd58908;
    data[13437] =  'sd79167;
    data[13438] =  'sd62646;
    data[13439] = -'sd53001;
    data[13440] = -'sd43325;
    data[13441] =  'sd24407;
    data[13442] =  'sd7008;
    data[13443] =  'sd49056;
    data[13444] =  'sd15710;
    data[13445] = -'sd53871;
    data[13446] = -'sd49415;
    data[13447] = -'sd18223;
    data[13448] =  'sd36280;
    data[13449] = -'sd73722;
    data[13450] = -'sd24531;
    data[13451] = -'sd7876;
    data[13452] = -'sd55132;
    data[13453] = -'sd58242;
    data[13454] = -'sd80012;
    data[13455] = -'sd68561;
    data[13456] =  'sd11596;
    data[13457] =  'sd81172;
    data[13458] =  'sd76681;
    data[13459] =  'sd45244;
    data[13460] = -'sd10974;
    data[13461] = -'sd76818;
    data[13462] = -'sd46203;
    data[13463] =  'sd4261;
    data[13464] =  'sd29827;
    data[13465] =  'sd44948;
    data[13466] = -'sd13046;
    data[13467] =  'sd72519;
    data[13468] =  'sd16110;
    data[13469] = -'sd51071;
    data[13470] = -'sd29815;
    data[13471] = -'sd44864;
    data[13472] =  'sd13634;
    data[13473] = -'sd68403;
    data[13474] =  'sd12702;
    data[13475] = -'sd74927;
    data[13476] = -'sd32966;
    data[13477] = -'sd66921;
    data[13478] =  'sd23076;
    data[13479] = -'sd2309;
    data[13480] = -'sd16163;
    data[13481] =  'sd50700;
    data[13482] =  'sd27218;
    data[13483] =  'sd26685;
    data[13484] =  'sd22954;
    data[13485] = -'sd3163;
    data[13486] = -'sd22141;
    data[13487] =  'sd8854;
    data[13488] =  'sd61978;
    data[13489] = -'sd57677;
    data[13490] = -'sd76057;
    data[13491] = -'sd40876;
    data[13492] =  'sd41550;
    data[13493] = -'sd36832;
    data[13494] =  'sd69858;
    data[13495] = -'sd2517;
    data[13496] = -'sd17619;
    data[13497] =  'sd40508;
    data[13498] = -'sd44126;
    data[13499] =  'sd18800;
    data[13500] = -'sd32241;
    data[13501] = -'sd61846;
    data[13502] =  'sd58601;
    data[13503] = -'sd81316;
    data[13504] = -'sd77689;
    data[13505] = -'sd52300;
    data[13506] = -'sd38418;
    data[13507] =  'sd58756;
    data[13508] = -'sd80231;
    data[13509] = -'sd70094;
    data[13510] =  'sd865;
    data[13511] =  'sd6055;
    data[13512] =  'sd42385;
    data[13513] = -'sd30987;
    data[13514] = -'sd53068;
    data[13515] = -'sd43794;
    data[13516] =  'sd21124;
    data[13517] = -'sd15973;
    data[13518] =  'sd52030;
    data[13519] =  'sd36528;
    data[13520] = -'sd71986;
    data[13521] = -'sd12379;
    data[13522] =  'sd77188;
    data[13523] =  'sd48793;
    data[13524] =  'sd13869;
    data[13525] = -'sd66758;
    data[13526] =  'sd24217;
    data[13527] =  'sd5678;
    data[13528] =  'sd39746;
    data[13529] = -'sd49460;
    data[13530] = -'sd18538;
    data[13531] =  'sd34075;
    data[13532] =  'sd74684;
    data[13533] =  'sd31265;
    data[13534] =  'sd55014;
    data[13535] =  'sd57416;
    data[13536] =  'sd74230;
    data[13537] =  'sd28087;
    data[13538] =  'sd32768;
    data[13539] =  'sd65535;
    data[13540] = -'sd32778;
    data[13541] = -'sd65605;
    data[13542] =  'sd32288;
    data[13543] =  'sd62175;
    data[13544] = -'sd56298;
    data[13545] = -'sd66404;
    data[13546] =  'sd26695;
    data[13547] =  'sd23024;
    data[13548] = -'sd2673;
    data[13549] = -'sd18711;
    data[13550] =  'sd32864;
    data[13551] =  'sd66207;
    data[13552] = -'sd28074;
    data[13553] = -'sd32677;
    data[13554] = -'sd64898;
    data[13555] =  'sd37237;
    data[13556] = -'sd67023;
    data[13557] =  'sd22362;
    data[13558] = -'sd7307;
    data[13559] = -'sd51149;
    data[13560] = -'sd30361;
    data[13561] = -'sd48686;
    data[13562] = -'sd13120;
    data[13563] =  'sd72001;
    data[13564] =  'sd12484;
    data[13565] = -'sd76453;
    data[13566] = -'sd43648;
    data[13567] =  'sd22146;
    data[13568] = -'sd8819;
    data[13569] = -'sd61733;
    data[13570] =  'sd59392;
    data[13571] = -'sd75779;
    data[13572] = -'sd38930;
    data[13573] =  'sd55172;
    data[13574] =  'sd58522;
    data[13575] = -'sd81869;
    data[13576] = -'sd81560;
    data[13577] = -'sd79397;
    data[13578] = -'sd64256;
    data[13579] =  'sd41731;
    data[13580] = -'sd35565;
    data[13581] =  'sd78727;
    data[13582] =  'sd59566;
    data[13583] = -'sd74561;
    data[13584] = -'sd30404;
    data[13585] = -'sd48987;
    data[13586] = -'sd15227;
    data[13587] =  'sd57252;
    data[13588] =  'sd73082;
    data[13589] =  'sd20051;
    data[13590] = -'sd23484;
    data[13591] = -'sd547;
    data[13592] = -'sd3829;
    data[13593] = -'sd26803;
    data[13594] = -'sd23780;
    data[13595] = -'sd2619;
    data[13596] = -'sd18333;
    data[13597] =  'sd35510;
    data[13598] = -'sd79112;
    data[13599] = -'sd62261;
    data[13600] =  'sd55696;
    data[13601] =  'sd62190;
    data[13602] = -'sd56193;
    data[13603] = -'sd65669;
    data[13604] =  'sd31840;
    data[13605] =  'sd59039;
    data[13606] = -'sd78250;
    data[13607] = -'sd56227;
    data[13608] = -'sd65907;
    data[13609] =  'sd30174;
    data[13610] =  'sd47377;
    data[13611] =  'sd3957;
    data[13612] =  'sd27699;
    data[13613] =  'sd30052;
    data[13614] =  'sd46523;
    data[13615] = -'sd2021;
    data[13616] = -'sd14147;
    data[13617] =  'sd64812;
    data[13618] = -'sd37839;
    data[13619] =  'sd62809;
    data[13620] = -'sd51860;
    data[13621] = -'sd35338;
    data[13622] =  'sd80316;
    data[13623] =  'sd70689;
    data[13624] =  'sd3300;
    data[13625] =  'sd23100;
    data[13626] = -'sd2141;
    data[13627] = -'sd14987;
    data[13628] =  'sd58932;
    data[13629] = -'sd78999;
    data[13630] = -'sd61470;
    data[13631] =  'sd61233;
    data[13632] = -'sd62892;
    data[13633] =  'sd51279;
    data[13634] =  'sd31271;
    data[13635] =  'sd55056;
    data[13636] =  'sd57710;
    data[13637] =  'sd76288;
    data[13638] =  'sd42493;
    data[13639] = -'sd30231;
    data[13640] = -'sd47776;
    data[13641] = -'sd6750;
    data[13642] = -'sd47250;
    data[13643] = -'sd3068;
    data[13644] = -'sd21476;
    data[13645] =  'sd13509;
    data[13646] = -'sd69278;
    data[13647] =  'sd6577;
    data[13648] =  'sd46039;
    data[13649] = -'sd5409;
    data[13650] = -'sd37863;
    data[13651] =  'sd62641;
    data[13652] = -'sd53036;
    data[13653] = -'sd43570;
    data[13654] =  'sd22692;
    data[13655] = -'sd4997;
    data[13656] = -'sd34979;
    data[13657] = -'sd81012;
    data[13658] = -'sd75561;
    data[13659] = -'sd37404;
    data[13660] =  'sd65854;
    data[13661] = -'sd30545;
    data[13662] = -'sd49974;
    data[13663] = -'sd22136;
    data[13664] =  'sd8889;
    data[13665] =  'sd62223;
    data[13666] = -'sd55962;
    data[13667] = -'sd64052;
    data[13668] =  'sd43159;
    data[13669] = -'sd25569;
    data[13670] = -'sd15142;
    data[13671] =  'sd57847;
    data[13672] =  'sd77247;
    data[13673] =  'sd49206;
    data[13674] =  'sd16760;
    data[13675] = -'sd46521;
    data[13676] =  'sd2035;
    data[13677] =  'sd14245;
    data[13678] = -'sd64126;
    data[13679] =  'sd42641;
    data[13680] = -'sd29195;
    data[13681] = -'sd40524;
    data[13682] =  'sd44014;
    data[13683] = -'sd19584;
    data[13684] =  'sd26753;
    data[13685] =  'sd23430;
    data[13686] =  'sd169;
    data[13687] =  'sd1183;
    data[13688] =  'sd8281;
    data[13689] =  'sd57967;
    data[13690] =  'sd78087;
    data[13691] =  'sd55086;
    data[13692] =  'sd57920;
    data[13693] =  'sd77758;
    data[13694] =  'sd52783;
    data[13695] =  'sd41799;
    data[13696] = -'sd35089;
    data[13697] = -'sd81782;
    data[13698] = -'sd80951;
    data[13699] = -'sd75134;
    data[13700] = -'sd34415;
    data[13701] = -'sd77064;
    data[13702] = -'sd47925;
    data[13703] = -'sd7793;
    data[13704] = -'sd54551;
    data[13705] = -'sd54175;
    data[13706] = -'sd51543;
    data[13707] = -'sd33119;
    data[13708] = -'sd67992;
    data[13709] =  'sd15579;
    data[13710] = -'sd54788;
    data[13711] = -'sd55834;
    data[13712] = -'sd63156;
    data[13713] =  'sd49431;
    data[13714] =  'sd18335;
    data[13715] = -'sd35496;
    data[13716] =  'sd79210;
    data[13717] =  'sd62947;
    data[13718] = -'sd50894;
    data[13719] = -'sd28576;
    data[13720] = -'sd36191;
    data[13721] =  'sd74345;
    data[13722] =  'sd28892;
    data[13723] =  'sd38403;
    data[13724] = -'sd58861;
    data[13725] =  'sd79496;
    data[13726] =  'sd64949;
    data[13727] = -'sd36880;
    data[13728] =  'sd69522;
    data[13729] = -'sd4869;
    data[13730] = -'sd34083;
    data[13731] = -'sd74740;
    data[13732] = -'sd31657;
    data[13733] = -'sd57758;
    data[13734] = -'sd76624;
    data[13735] = -'sd44845;
    data[13736] =  'sd13767;
    data[13737] = -'sd67472;
    data[13738] =  'sd19219;
    data[13739] = -'sd29308;
    data[13740] = -'sd41315;
    data[13741] =  'sd38477;
    data[13742] = -'sd58343;
    data[13743] = -'sd80719;
    data[13744] = -'sd73510;
    data[13745] = -'sd23047;
    data[13746] =  'sd2512;
    data[13747] =  'sd17584;
    data[13748] = -'sd40753;
    data[13749] =  'sd42411;
    data[13750] = -'sd30805;
    data[13751] = -'sd51794;
    data[13752] = -'sd34876;
    data[13753] = -'sd80291;
    data[13754] = -'sd70514;
    data[13755] = -'sd2075;
    data[13756] = -'sd14525;
    data[13757] =  'sd62166;
    data[13758] = -'sd56361;
    data[13759] = -'sd66845;
    data[13760] =  'sd23608;
    data[13761] =  'sd1415;
    data[13762] =  'sd9905;
    data[13763] =  'sd69335;
    data[13764] = -'sd6178;
    data[13765] = -'sd43246;
    data[13766] =  'sd24960;
    data[13767] =  'sd10879;
    data[13768] =  'sd76153;
    data[13769] =  'sd41548;
    data[13770] = -'sd36846;
    data[13771] =  'sd69760;
    data[13772] = -'sd3203;
    data[13773] = -'sd22421;
    data[13774] =  'sd6894;
    data[13775] =  'sd48258;
    data[13776] =  'sd10124;
    data[13777] =  'sd70868;
    data[13778] =  'sd4553;
    data[13779] =  'sd31871;
    data[13780] =  'sd59256;
    data[13781] = -'sd76731;
    data[13782] = -'sd45594;
    data[13783] =  'sd8524;
    data[13784] =  'sd59668;
    data[13785] = -'sd73847;
    data[13786] = -'sd25406;
    data[13787] = -'sd14001;
    data[13788] =  'sd65834;
    data[13789] = -'sd30685;
    data[13790] = -'sd50954;
    data[13791] = -'sd28996;
    data[13792] = -'sd39131;
    data[13793] =  'sd53765;
    data[13794] =  'sd48673;
    data[13795] =  'sd13029;
    data[13796] = -'sd72638;
    data[13797] = -'sd16943;
    data[13798] =  'sd45240;
    data[13799] = -'sd11002;
    data[13800] = -'sd77014;
    data[13801] = -'sd47575;
    data[13802] = -'sd5343;
    data[13803] = -'sd37401;
    data[13804] =  'sd65875;
    data[13805] = -'sd30398;
    data[13806] = -'sd48945;
    data[13807] = -'sd14933;
    data[13808] =  'sd59310;
    data[13809] = -'sd76353;
    data[13810] = -'sd42948;
    data[13811] =  'sd27046;
    data[13812] =  'sd25481;
    data[13813] =  'sd14526;
    data[13814] = -'sd62159;
    data[13815] =  'sd56410;
    data[13816] =  'sd67188;
    data[13817] = -'sd21207;
    data[13818] =  'sd15392;
    data[13819] = -'sd56097;
    data[13820] = -'sd64997;
    data[13821] =  'sd36544;
    data[13822] = -'sd71874;
    data[13823] = -'sd11595;
    data[13824] = -'sd81165;
    data[13825] = -'sd76632;
    data[13826] = -'sd44901;
    data[13827] =  'sd13375;
    data[13828] = -'sd70216;
    data[13829] =  'sd11;
    data[13830] =  'sd77;
    data[13831] =  'sd539;
    data[13832] =  'sd3773;
    data[13833] =  'sd26411;
    data[13834] =  'sd21036;
    data[13835] = -'sd16589;
    data[13836] =  'sd47718;
    data[13837] =  'sd6344;
    data[13838] =  'sd44408;
    data[13839] = -'sd16826;
    data[13840] =  'sd46059;
    data[13841] = -'sd5269;
    data[13842] = -'sd36883;
    data[13843] =  'sd69501;
    data[13844] = -'sd5016;
    data[13845] = -'sd35112;
    data[13846] =  'sd81898;
    data[13847] =  'sd81763;
    data[13848] =  'sd80818;
    data[13849] =  'sd74203;
    data[13850] =  'sd27898;
    data[13851] =  'sd31445;
    data[13852] =  'sd56274;
    data[13853] =  'sd66236;
    data[13854] = -'sd27871;
    data[13855] = -'sd31256;
    data[13856] = -'sd54951;
    data[13857] = -'sd56975;
    data[13858] = -'sd71143;
    data[13859] = -'sd6478;
    data[13860] = -'sd45346;
    data[13861] =  'sd10260;
    data[13862] =  'sd71820;
    data[13863] =  'sd11217;
    data[13864] =  'sd78519;
    data[13865] =  'sd58110;
    data[13866] =  'sd79088;
    data[13867] =  'sd62093;
    data[13868] = -'sd56872;
    data[13869] = -'sd70422;
    data[13870] = -'sd1431;
    data[13871] = -'sd10017;
    data[13872] = -'sd70119;
    data[13873] =  'sd690;
    data[13874] =  'sd4830;
    data[13875] =  'sd33810;
    data[13876] =  'sd72829;
    data[13877] =  'sd18280;
    data[13878] = -'sd35881;
    data[13879] =  'sd76515;
    data[13880] =  'sd44082;
    data[13881] = -'sd19108;
    data[13882] =  'sd30085;
    data[13883] =  'sd46754;
    data[13884] = -'sd404;
    data[13885] = -'sd2828;
    data[13886] = -'sd19796;
    data[13887] =  'sd25269;
    data[13888] =  'sd13042;
    data[13889] = -'sd72547;
    data[13890] = -'sd16306;
    data[13891] =  'sd49699;
    data[13892] =  'sd20211;
    data[13893] = -'sd22364;
    data[13894] =  'sd7293;
    data[13895] =  'sd51051;
    data[13896] =  'sd29675;
    data[13897] =  'sd43884;
    data[13898] = -'sd20494;
    data[13899] =  'sd20383;
    data[13900] = -'sd21160;
    data[13901] =  'sd15721;
    data[13902] = -'sd53794;
    data[13903] = -'sd48876;
    data[13904] = -'sd14450;
    data[13905] =  'sd62691;
    data[13906] = -'sd52686;
    data[13907] = -'sd41120;
    data[13908] =  'sd39842;
    data[13909] = -'sd48788;
    data[13910] = -'sd13834;
    data[13911] =  'sd67003;
    data[13912] = -'sd22502;
    data[13913] =  'sd6327;
    data[13914] =  'sd44289;
    data[13915] = -'sd17659;
    data[13916] =  'sd40228;
    data[13917] = -'sd46086;
    data[13918] =  'sd5080;
    data[13919] =  'sd35560;
    data[13920] = -'sd78762;
    data[13921] = -'sd59811;
    data[13922] =  'sd72846;
    data[13923] =  'sd18399;
    data[13924] = -'sd35048;
    data[13925] = -'sd81495;
    data[13926] = -'sd78942;
    data[13927] = -'sd61071;
    data[13928] =  'sd64026;
    data[13929] = -'sd43341;
    data[13930] =  'sd24295;
    data[13931] =  'sd6224;
    data[13932] =  'sd43568;
    data[13933] = -'sd22706;
    data[13934] =  'sd4899;
    data[13935] =  'sd34293;
    data[13936] =  'sd76210;
    data[13937] =  'sd41947;
    data[13938] = -'sd34053;
    data[13939] = -'sd74530;
    data[13940] = -'sd30187;
    data[13941] = -'sd47468;
    data[13942] = -'sd4594;
    data[13943] = -'sd32158;
    data[13944] = -'sd61265;
    data[13945] =  'sd62668;
    data[13946] = -'sd52847;
    data[13947] = -'sd42247;
    data[13948] =  'sd31953;
    data[13949] =  'sd59830;
    data[13950] = -'sd72713;
    data[13951] = -'sd17468;
    data[13952] =  'sd41565;
    data[13953] = -'sd36727;
    data[13954] =  'sd70593;
    data[13955] =  'sd2628;
    data[13956] =  'sd18396;
    data[13957] = -'sd35069;
    data[13958] = -'sd81642;
    data[13959] = -'sd79971;
    data[13960] = -'sd68274;
    data[13961] =  'sd13605;
    data[13962] = -'sd68606;
    data[13963] =  'sd11281;
    data[13964] =  'sd78967;
    data[13965] =  'sd61246;
    data[13966] = -'sd62801;
    data[13967] =  'sd51916;
    data[13968] =  'sd35730;
    data[13969] = -'sd77572;
    data[13970] = -'sd51481;
    data[13971] = -'sd32685;
    data[13972] = -'sd64954;
    data[13973] =  'sd36845;
    data[13974] = -'sd69767;
    data[13975] =  'sd3154;
    data[13976] =  'sd22078;
    data[13977] = -'sd9295;
    data[13978] = -'sd65065;
    data[13979] =  'sd36068;
    data[13980] = -'sd75206;
    data[13981] = -'sd34919;
    data[13982] = -'sd80592;
    data[13983] = -'sd72621;
    data[13984] = -'sd16824;
    data[13985] =  'sd46073;
    data[13986] = -'sd5171;
    data[13987] = -'sd36197;
    data[13988] =  'sd74303;
    data[13989] =  'sd28598;
    data[13990] =  'sd36345;
    data[13991] = -'sd73267;
    data[13992] = -'sd21346;
    data[13993] =  'sd14419;
    data[13994] = -'sd62908;
    data[13995] =  'sd51167;
    data[13996] =  'sd30487;
    data[13997] =  'sd49568;
    data[13998] =  'sd19294;
    data[13999] = -'sd28783;
    data[14000] = -'sd37640;
    data[14001] =  'sd64202;
    data[14002] = -'sd42109;
    data[14003] =  'sd32919;
    data[14004] =  'sd66592;
    data[14005] = -'sd25379;
    data[14006] = -'sd13812;
    data[14007] =  'sd67157;
    data[14008] = -'sd21424;
    data[14009] =  'sd13873;
    data[14010] = -'sd66730;
    data[14011] =  'sd24413;
    data[14012] =  'sd7050;
    data[14013] =  'sd49350;
    data[14014] =  'sd17768;
    data[14015] = -'sd39465;
    data[14016] =  'sd51427;
    data[14017] =  'sd32307;
    data[14018] =  'sd62308;
    data[14019] = -'sd55367;
    data[14020] = -'sd59887;
    data[14021] =  'sd72314;
    data[14022] =  'sd14675;
    data[14023] = -'sd61116;
    data[14024] =  'sd63711;
    data[14025] = -'sd45546;
    data[14026] =  'sd8860;
    data[14027] =  'sd62020;
    data[14028] = -'sd57383;
    data[14029] = -'sd73999;
    data[14030] = -'sd26470;
    data[14031] = -'sd21449;
    data[14032] =  'sd13698;
    data[14033] = -'sd67955;
    data[14034] =  'sd15838;
    data[14035] = -'sd52975;
    data[14036] = -'sd43143;
    data[14037] =  'sd25681;
    data[14038] =  'sd15926;
    data[14039] = -'sd52359;
    data[14040] = -'sd38831;
    data[14041] =  'sd55865;
    data[14042] =  'sd63373;
    data[14043] = -'sd47912;
    data[14044] = -'sd7702;
    data[14045] = -'sd53914;
    data[14046] = -'sd49716;
    data[14047] = -'sd20330;
    data[14048] =  'sd21531;
    data[14049] = -'sd13124;
    data[14050] =  'sd71973;
    data[14051] =  'sd12288;
    data[14052] = -'sd77825;
    data[14053] = -'sd53252;
    data[14054] = -'sd45082;
    data[14055] =  'sd12108;
    data[14056] = -'sd79085;
    data[14057] = -'sd62072;
    data[14058] =  'sd57019;
    data[14059] =  'sd71451;
    data[14060] =  'sd8634;
    data[14061] =  'sd60438;
    data[14062] = -'sd68457;
    data[14063] =  'sd12324;
    data[14064] = -'sd77573;
    data[14065] = -'sd51488;
    data[14066] = -'sd32734;
    data[14067] = -'sd65297;
    data[14068] =  'sd34444;
    data[14069] =  'sd77267;
    data[14070] =  'sd49346;
    data[14071] =  'sd17740;
    data[14072] = -'sd39661;
    data[14073] =  'sd50055;
    data[14074] =  'sd22703;
    data[14075] = -'sd4920;
    data[14076] = -'sd34440;
    data[14077] = -'sd77239;
    data[14078] = -'sd49150;
    data[14079] = -'sd16368;
    data[14080] =  'sd49265;
    data[14081] =  'sd17173;
    data[14082] = -'sd43630;
    data[14083] =  'sd22272;
    data[14084] = -'sd7937;
    data[14085] = -'sd55559;
    data[14086] = -'sd61231;
    data[14087] =  'sd62906;
    data[14088] = -'sd51181;
    data[14089] = -'sd30585;
    data[14090] = -'sd50254;
    data[14091] = -'sd24096;
    data[14092] = -'sd4831;
    data[14093] = -'sd33817;
    data[14094] = -'sd72878;
    data[14095] = -'sd18623;
    data[14096] =  'sd33480;
    data[14097] =  'sd70519;
    data[14098] =  'sd2110;
    data[14099] =  'sd14770;
    data[14100] = -'sd60451;
    data[14101] =  'sd68366;
    data[14102] = -'sd12961;
    data[14103] =  'sd73114;
    data[14104] =  'sd20275;
    data[14105] = -'sd21916;
    data[14106] =  'sd10429;
    data[14107] =  'sd73003;
    data[14108] =  'sd19498;
    data[14109] = -'sd27355;
    data[14110] = -'sd27644;
    data[14111] = -'sd29667;
    data[14112] = -'sd43828;
    data[14113] =  'sd20886;
    data[14114] = -'sd17639;
    data[14115] =  'sd40368;
    data[14116] = -'sd45106;
    data[14117] =  'sd11940;
    data[14118] = -'sd80261;
    data[14119] = -'sd70304;
    data[14120] = -'sd605;
    data[14121] = -'sd4235;
    data[14122] = -'sd29645;
    data[14123] = -'sd43674;
    data[14124] =  'sd21964;
    data[14125] = -'sd10093;
    data[14126] = -'sd70651;
    data[14127] = -'sd3034;
    data[14128] = -'sd21238;
    data[14129] =  'sd15175;
    data[14130] = -'sd57616;
    data[14131] = -'sd75630;
    data[14132] = -'sd37887;
    data[14133] =  'sd62473;
    data[14134] = -'sd54212;
    data[14135] = -'sd51802;
    data[14136] = -'sd34932;
    data[14137] = -'sd80683;
    data[14138] = -'sd73258;
    data[14139] = -'sd21283;
    data[14140] =  'sd14860;
    data[14141] = -'sd59821;
    data[14142] =  'sd72776;
    data[14143] =  'sd17909;
    data[14144] = -'sd38478;
    data[14145] =  'sd58336;
    data[14146] =  'sd80670;
    data[14147] =  'sd73167;
    data[14148] =  'sd20646;
    data[14149] = -'sd19319;
    data[14150] =  'sd28608;
    data[14151] =  'sd36415;
    data[14152] = -'sd72777;
    data[14153] = -'sd17916;
    data[14154] =  'sd38429;
    data[14155] = -'sd58679;
    data[14156] =  'sd80770;
    data[14157] =  'sd73867;
    data[14158] =  'sd25546;
    data[14159] =  'sd14981;
    data[14160] = -'sd58974;
    data[14161] =  'sd78705;
    data[14162] =  'sd59412;
    data[14163] = -'sd75639;
    data[14164] = -'sd37950;
    data[14165] =  'sd62032;
    data[14166] = -'sd57299;
    data[14167] = -'sd73411;
    data[14168] = -'sd22354;
    data[14169] =  'sd7363;
    data[14170] =  'sd51541;
    data[14171] =  'sd33105;
    data[14172] =  'sd67894;
    data[14173] = -'sd16265;
    data[14174] =  'sd49986;
    data[14175] =  'sd22220;
    data[14176] = -'sd8301;
    data[14177] = -'sd58107;
    data[14178] = -'sd79067;
    data[14179] = -'sd61946;
    data[14180] =  'sd57901;
    data[14181] =  'sd77625;
    data[14182] =  'sd51852;
    data[14183] =  'sd35282;
    data[14184] = -'sd80708;
    data[14185] = -'sd73433;
    data[14186] = -'sd22508;
    data[14187] =  'sd6285;
    data[14188] =  'sd43995;
    data[14189] = -'sd19717;
    data[14190] =  'sd25822;
    data[14191] =  'sd16913;
    data[14192] = -'sd45450;
    data[14193] =  'sd9532;
    data[14194] =  'sd66724;
    data[14195] = -'sd24455;
    data[14196] = -'sd7344;
    data[14197] = -'sd51408;
    data[14198] = -'sd32174;
    data[14199] = -'sd61377;
    data[14200] =  'sd61884;
    data[14201] = -'sd58335;
    data[14202] = -'sd80663;
    data[14203] = -'sd73118;
    data[14204] = -'sd20303;
    data[14205] =  'sd21720;
    data[14206] = -'sd11801;
    data[14207] =  'sd81234;
    data[14208] =  'sd77115;
    data[14209] =  'sd48282;
    data[14210] =  'sd10292;
    data[14211] =  'sd72044;
    data[14212] =  'sd12785;
    data[14213] = -'sd74346;
    data[14214] = -'sd28899;
    data[14215] = -'sd38452;
    data[14216] =  'sd58518;
    data[14217] = -'sd81897;
    data[14218] = -'sd81756;
    data[14219] = -'sd80769;
    data[14220] = -'sd73860;
    data[14221] = -'sd25497;
    data[14222] = -'sd14638;
    data[14223] =  'sd61375;
    data[14224] = -'sd61898;
    data[14225] =  'sd58237;
    data[14226] =  'sd79977;
    data[14227] =  'sd68316;
    data[14228] = -'sd13311;
    data[14229] =  'sd70664;
    data[14230] =  'sd3125;
    data[14231] =  'sd21875;
    data[14232] = -'sd10716;
    data[14233] = -'sd75012;
    data[14234] = -'sd33561;
    data[14235] = -'sd71086;
    data[14236] = -'sd6079;
    data[14237] = -'sd42553;
    data[14238] =  'sd29811;
    data[14239] =  'sd44836;
    data[14240] = -'sd13830;
    data[14241] =  'sd67031;
    data[14242] = -'sd22306;
    data[14243] =  'sd7699;
    data[14244] =  'sd53893;
    data[14245] =  'sd49569;
    data[14246] =  'sd19301;
    data[14247] = -'sd28734;
    data[14248] = -'sd37297;
    data[14249] =  'sd66603;
    data[14250] = -'sd25302;
    data[14251] = -'sd13273;
    data[14252] =  'sd70930;
    data[14253] =  'sd4987;
    data[14254] =  'sd34909;
    data[14255] =  'sd80522;
    data[14256] =  'sd72131;
    data[14257] =  'sd13394;
    data[14258] = -'sd70083;
    data[14259] =  'sd942;
    data[14260] =  'sd6594;
    data[14261] =  'sd46158;
    data[14262] = -'sd4576;
    data[14263] = -'sd32032;
    data[14264] = -'sd60383;
    data[14265] =  'sd68842;
    data[14266] = -'sd9629;
    data[14267] = -'sd67403;
    data[14268] =  'sd19702;
    data[14269] = -'sd25927;
    data[14270] = -'sd17648;
    data[14271] =  'sd40305;
    data[14272] = -'sd45547;
    data[14273] =  'sd8853;
    data[14274] =  'sd61971;
    data[14275] = -'sd57726;
    data[14276] = -'sd76400;
    data[14277] = -'sd43277;
    data[14278] =  'sd24743;
    data[14279] =  'sd9360;
    data[14280] =  'sd65520;
    data[14281] = -'sd32883;
    data[14282] = -'sd66340;
    data[14283] =  'sd27143;
    data[14284] =  'sd26160;
    data[14285] =  'sd19279;
    data[14286] = -'sd28888;
    data[14287] = -'sd38375;
    data[14288] =  'sd59057;
    data[14289] = -'sd78124;
    data[14290] = -'sd55345;
    data[14291] = -'sd59733;
    data[14292] =  'sd73392;
    data[14293] =  'sd22221;
    data[14294] = -'sd8294;
    data[14295] = -'sd58058;
    data[14296] = -'sd78724;
    data[14297] = -'sd59545;
    data[14298] =  'sd74708;
    data[14299] =  'sd31433;
    data[14300] =  'sd56190;
    data[14301] =  'sd65648;
    data[14302] = -'sd31987;
    data[14303] = -'sd60068;
    data[14304] =  'sd71047;
    data[14305] =  'sd5806;
    data[14306] =  'sd40642;
    data[14307] = -'sd43188;
    data[14308] =  'sd25366;
    data[14309] =  'sd13721;
    data[14310] = -'sd67794;
    data[14311] =  'sd16965;
    data[14312] = -'sd45086;
    data[14313] =  'sd12080;
    data[14314] = -'sd79281;
    data[14315] = -'sd63444;
    data[14316] =  'sd47415;
    data[14317] =  'sd4223;
    data[14318] =  'sd29561;
    data[14319] =  'sd43086;
    data[14320] = -'sd26080;
    data[14321] = -'sd18719;
    data[14322] =  'sd32808;
    data[14323] =  'sd65815;
    data[14324] = -'sd30818;
    data[14325] = -'sd51885;
    data[14326] = -'sd35513;
    data[14327] =  'sd79091;
    data[14328] =  'sd62114;
    data[14329] = -'sd56725;
    data[14330] = -'sd69393;
    data[14331] =  'sd5772;
    data[14332] =  'sd40404;
    data[14333] = -'sd44854;
    data[14334] =  'sd13704;
    data[14335] = -'sd67913;
    data[14336] =  'sd16132;
    data[14337] = -'sd50917;
    data[14338] = -'sd28737;
    data[14339] = -'sd37318;
    data[14340] =  'sd66456;
    data[14341] = -'sd26331;
    data[14342] = -'sd20476;
    data[14343] =  'sd20509;
    data[14344] = -'sd20278;
    data[14345] =  'sd21895;
    data[14346] = -'sd10576;
    data[14347] = -'sd74032;
    data[14348] = -'sd26701;
    data[14349] = -'sd23066;
    data[14350] =  'sd2379;
    data[14351] =  'sd16653;
    data[14352] = -'sd47270;
    data[14353] = -'sd3208;
    data[14354] = -'sd22456;
    data[14355] =  'sd6649;
    data[14356] =  'sd46543;
    data[14357] = -'sd1881;
    data[14358] = -'sd13167;
    data[14359] =  'sd71672;
    data[14360] =  'sd10181;
    data[14361] =  'sd71267;
    data[14362] =  'sd7346;
    data[14363] =  'sd51422;
    data[14364] =  'sd32272;
    data[14365] =  'sd62063;
    data[14366] = -'sd57082;
    data[14367] = -'sd71892;
    data[14368] = -'sd11721;
    data[14369] =  'sd81794;
    data[14370] =  'sd81035;
    data[14371] =  'sd75722;
    data[14372] =  'sd38531;
    data[14373] = -'sd57965;
    data[14374] = -'sd78073;
    data[14375] = -'sd54988;
    data[14376] = -'sd57234;
    data[14377] = -'sd72956;
    data[14378] = -'sd19169;
    data[14379] =  'sd29658;
    data[14380] =  'sd43765;
    data[14381] = -'sd21327;
    data[14382] =  'sd14552;
    data[14383] = -'sd61977;
    data[14384] =  'sd57684;
    data[14385] =  'sd76106;
    data[14386] =  'sd41219;
    data[14387] = -'sd39149;
    data[14388] =  'sd53639;
    data[14389] =  'sd47791;
    data[14390] =  'sd6855;
    data[14391] =  'sd47985;
    data[14392] =  'sd8213;
    data[14393] =  'sd57491;
    data[14394] =  'sd74755;
    data[14395] =  'sd31762;
    data[14396] =  'sd58493;
    data[14397] =  'sd81769;
    data[14398] =  'sd80860;
    data[14399] =  'sd74497;
    data[14400] =  'sd29956;
    data[14401] =  'sd45851;
    data[14402] = -'sd6725;
    data[14403] = -'sd47075;
    data[14404] = -'sd1843;
    data[14405] = -'sd12901;
    data[14406] =  'sd73534;
    data[14407] =  'sd23215;
    data[14408] = -'sd1336;
    data[14409] = -'sd9352;
    data[14410] = -'sd65464;
    data[14411] =  'sd33275;
    data[14412] =  'sd69084;
    data[14413] = -'sd7935;
    data[14414] = -'sd55545;
    data[14415] = -'sd61133;
    data[14416] =  'sd63592;
    data[14417] = -'sd46379;
    data[14418] =  'sd3029;
    data[14419] =  'sd21203;
    data[14420] = -'sd15420;
    data[14421] =  'sd55901;
    data[14422] =  'sd63625;
    data[14423] = -'sd46148;
    data[14424] =  'sd4646;
    data[14425] =  'sd32522;
    data[14426] =  'sd63813;
    data[14427] = -'sd44832;
    data[14428] =  'sd13858;
    data[14429] = -'sd66835;
    data[14430] =  'sd23678;
    data[14431] =  'sd1905;
    data[14432] =  'sd13335;
    data[14433] = -'sd70496;
    data[14434] = -'sd1949;
    data[14435] = -'sd13643;
    data[14436] =  'sd68340;
    data[14437] = -'sd13143;
    data[14438] =  'sd71840;
    data[14439] =  'sd11357;
    data[14440] =  'sd79499;
    data[14441] =  'sd64970;
    data[14442] = -'sd36733;
    data[14443] =  'sd70551;
    data[14444] =  'sd2334;
    data[14445] =  'sd16338;
    data[14446] = -'sd49475;
    data[14447] = -'sd18643;
    data[14448] =  'sd33340;
    data[14449] =  'sd69539;
    data[14450] = -'sd4750;
    data[14451] = -'sd33250;
    data[14452] = -'sd68909;
    data[14453] =  'sd9160;
    data[14454] =  'sd64120;
    data[14455] = -'sd42683;
    data[14456] =  'sd28901;
    data[14457] =  'sd38466;
    data[14458] = -'sd58420;
    data[14459] = -'sd81258;
    data[14460] = -'sd77283;
    data[14461] = -'sd49458;
    data[14462] = -'sd18524;
    data[14463] =  'sd34173;
    data[14464] =  'sd75370;
    data[14465] =  'sd36067;
    data[14466] = -'sd75213;
    data[14467] = -'sd34968;
    data[14468] = -'sd80935;
    data[14469] = -'sd75022;
    data[14470] = -'sd33631;
    data[14471] = -'sd71576;
    data[14472] = -'sd9509;
    data[14473] = -'sd66563;
    data[14474] =  'sd25582;
    data[14475] =  'sd15233;
    data[14476] = -'sd57210;
    data[14477] = -'sd72788;
    data[14478] = -'sd17993;
    data[14479] =  'sd37890;
    data[14480] = -'sd62452;
    data[14481] =  'sd54359;
    data[14482] =  'sd52831;
    data[14483] =  'sd42135;
    data[14484] = -'sd32737;
    data[14485] = -'sd65318;
    data[14486] =  'sd34297;
    data[14487] =  'sd76238;
    data[14488] =  'sd42143;
    data[14489] = -'sd32681;
    data[14490] = -'sd64926;
    data[14491] =  'sd37041;
    data[14492] = -'sd68395;
    data[14493] =  'sd12758;
    data[14494] = -'sd74535;
    data[14495] = -'sd30222;
    data[14496] = -'sd47713;
    data[14497] = -'sd6309;
    data[14498] = -'sd44163;
    data[14499] =  'sd18541;
    data[14500] = -'sd34054;
    data[14501] = -'sd74537;
    data[14502] = -'sd30236;
    data[14503] = -'sd47811;
    data[14504] = -'sd6995;
    data[14505] = -'sd48965;
    data[14506] = -'sd15073;
    data[14507] =  'sd58330;
    data[14508] =  'sd80628;
    data[14509] =  'sd72873;
    data[14510] =  'sd18588;
    data[14511] = -'sd33725;
    data[14512] = -'sd72234;
    data[14513] = -'sd14115;
    data[14514] =  'sd65036;
    data[14515] = -'sd36271;
    data[14516] =  'sd73785;
    data[14517] =  'sd24972;
    data[14518] =  'sd10963;
    data[14519] =  'sd76741;
    data[14520] =  'sd45664;
    data[14521] = -'sd8034;
    data[14522] = -'sd56238;
    data[14523] = -'sd65984;
    data[14524] =  'sd29635;
    data[14525] =  'sd43604;
    data[14526] = -'sd22454;
    data[14527] =  'sd6663;
    data[14528] =  'sd46641;
    data[14529] = -'sd1195;
    data[14530] = -'sd8365;
    data[14531] = -'sd58555;
    data[14532] =  'sd81638;
    data[14533] =  'sd79943;
    data[14534] =  'sd68078;
    data[14535] = -'sd14977;
    data[14536] =  'sd59002;
    data[14537] = -'sd78509;
    data[14538] = -'sd58040;
    data[14539] = -'sd78598;
    data[14540] = -'sd58663;
    data[14541] =  'sd80882;
    data[14542] =  'sd74651;
    data[14543] =  'sd31034;
    data[14544] =  'sd53397;
    data[14545] =  'sd46097;
    data[14546] = -'sd5003;
    data[14547] = -'sd35021;
    data[14548] = -'sd81306;
    data[14549] = -'sd77619;
    data[14550] = -'sd51810;
    data[14551] = -'sd34988;
    data[14552] = -'sd81075;
    data[14553] = -'sd76002;
    data[14554] = -'sd40491;
    data[14555] =  'sd44245;
    data[14556] = -'sd17967;
    data[14557] =  'sd38072;
    data[14558] = -'sd61178;
    data[14559] =  'sd63277;
    data[14560] = -'sd48584;
    data[14561] = -'sd12406;
    data[14562] =  'sd76999;
    data[14563] =  'sd47470;
    data[14564] =  'sd4608;
    data[14565] =  'sd32256;
    data[14566] =  'sd61951;
    data[14567] = -'sd57866;
    data[14568] = -'sd77380;
    data[14569] = -'sd50137;
    data[14570] = -'sd23277;
    data[14571] =  'sd902;
    data[14572] =  'sd6314;
    data[14573] =  'sd44198;
    data[14574] = -'sd18296;
    data[14575] =  'sd35769;
    data[14576] = -'sd77299;
    data[14577] = -'sd49570;
    data[14578] = -'sd19308;
    data[14579] =  'sd28685;
    data[14580] =  'sd36954;
    data[14581] = -'sd69004;
    data[14582] =  'sd8495;
    data[14583] =  'sd59465;
    data[14584] = -'sd75268;
    data[14585] = -'sd35353;
    data[14586] =  'sd80211;
    data[14587] =  'sd69954;
    data[14588] = -'sd1845;
    data[14589] = -'sd12915;
    data[14590] =  'sd73436;
    data[14591] =  'sd22529;
    data[14592] = -'sd6138;
    data[14593] = -'sd42966;
    data[14594] =  'sd26920;
    data[14595] =  'sd24599;
    data[14596] =  'sd8352;
    data[14597] =  'sd58464;
    data[14598] =  'sd81566;
    data[14599] =  'sd79439;
    data[14600] =  'sd64550;
    data[14601] = -'sd39673;
    data[14602] =  'sd49971;
    data[14603] =  'sd22115;
    data[14604] = -'sd9036;
    data[14605] = -'sd63252;
    data[14606] =  'sd48759;
    data[14607] =  'sd13631;
    data[14608] = -'sd68424;
    data[14609] =  'sd12555;
    data[14610] = -'sd75956;
    data[14611] = -'sd40169;
    data[14612] =  'sd46499;
    data[14613] = -'sd2189;
    data[14614] = -'sd15323;
    data[14615] =  'sd56580;
    data[14616] =  'sd68378;
    data[14617] = -'sd12877;
    data[14618] =  'sd73702;
    data[14619] =  'sd24391;
    data[14620] =  'sd6896;
    data[14621] =  'sd48272;
    data[14622] =  'sd10222;
    data[14623] =  'sd71554;
    data[14624] =  'sd9355;
    data[14625] =  'sd65485;
    data[14626] = -'sd33128;
    data[14627] = -'sd68055;
    data[14628] =  'sd15138;
    data[14629] = -'sd57875;
    data[14630] = -'sd77443;
    data[14631] = -'sd50578;
    data[14632] = -'sd26364;
    data[14633] = -'sd20707;
    data[14634] =  'sd18892;
    data[14635] = -'sd31597;
    data[14636] = -'sd57338;
    data[14637] = -'sd73684;
    data[14638] = -'sd24265;
    data[14639] = -'sd6014;
    data[14640] = -'sd42098;
    data[14641] =  'sd32996;
    data[14642] =  'sd67131;
    data[14643] = -'sd21606;
    data[14644] =  'sd12599;
    data[14645] = -'sd75648;
    data[14646] = -'sd38013;
    data[14647] =  'sd61591;
    data[14648] = -'sd60386;
    data[14649] =  'sd68821;
    data[14650] = -'sd9776;
    data[14651] = -'sd68432;
    data[14652] =  'sd12499;
    data[14653] = -'sd76348;
    data[14654] = -'sd42913;
    data[14655] =  'sd27291;
    data[14656] =  'sd27196;
    data[14657] =  'sd26531;
    data[14658] =  'sd21876;
    data[14659] = -'sd10709;
    data[14660] = -'sd74963;
    data[14661] = -'sd33218;
    data[14662] = -'sd68685;
    data[14663] =  'sd10728;
    data[14664] =  'sd75096;
    data[14665] =  'sd34149;
    data[14666] =  'sd75202;
    data[14667] =  'sd34891;
    data[14668] =  'sd80396;
    data[14669] =  'sd71249;
    data[14670] =  'sd7220;
    data[14671] =  'sd50540;
    data[14672] =  'sd26098;
    data[14673] =  'sd18845;
    data[14674] = -'sd31926;
    data[14675] = -'sd59641;
    data[14676] =  'sd74036;
    data[14677] =  'sd26729;
    data[14678] =  'sd23262;
    data[14679] = -'sd1007;
    data[14680] = -'sd7049;
    data[14681] = -'sd49343;
    data[14682] = -'sd17719;
    data[14683] =  'sd39808;
    data[14684] = -'sd49026;
    data[14685] = -'sd15500;
    data[14686] =  'sd55341;
    data[14687] =  'sd59705;
    data[14688] = -'sd73588;
    data[14689] = -'sd23593;
    data[14690] = -'sd1310;
    data[14691] = -'sd9170;
    data[14692] = -'sd64190;
    data[14693] =  'sd42193;
    data[14694] = -'sd32331;
    data[14695] = -'sd62476;
    data[14696] =  'sd54191;
    data[14697] =  'sd51655;
    data[14698] =  'sd33903;
    data[14699] =  'sd73480;
    data[14700] =  'sd22837;
    data[14701] = -'sd3982;
    data[14702] = -'sd27874;
    data[14703] = -'sd31277;
    data[14704] = -'sd55098;
    data[14705] = -'sd58004;
    data[14706] = -'sd78346;
    data[14707] = -'sd56899;
    data[14708] = -'sd70611;
    data[14709] = -'sd2754;
    data[14710] = -'sd19278;
    data[14711] =  'sd28895;
    data[14712] =  'sd38424;
    data[14713] = -'sd58714;
    data[14714] =  'sd80525;
    data[14715] =  'sd72152;
    data[14716] =  'sd13541;
    data[14717] = -'sd69054;
    data[14718] =  'sd8145;
    data[14719] =  'sd57015;
    data[14720] =  'sd71423;
    data[14721] =  'sd8438;
    data[14722] =  'sd59066;
    data[14723] = -'sd78061;
    data[14724] = -'sd54904;
    data[14725] = -'sd56646;
    data[14726] = -'sd68840;
    data[14727] =  'sd9643;
    data[14728] =  'sd67501;
    data[14729] = -'sd19016;
    data[14730] =  'sd30729;
    data[14731] =  'sd51262;
    data[14732] =  'sd31152;
    data[14733] =  'sd54223;
    data[14734] =  'sd51879;
    data[14735] =  'sd35471;
    data[14736] = -'sd79385;
    data[14737] = -'sd64172;
    data[14738] =  'sd42319;
    data[14739] = -'sd31449;
    data[14740] = -'sd56302;
    data[14741] = -'sd66432;
    data[14742] =  'sd26499;
    data[14743] =  'sd21652;
    data[14744] = -'sd12277;
    data[14745] =  'sd77902;
    data[14746] =  'sd53791;
    data[14747] =  'sd48855;
    data[14748] =  'sd14303;
    data[14749] = -'sd63720;
    data[14750] =  'sd45483;
    data[14751] = -'sd9301;
    data[14752] = -'sd65107;
    data[14753] =  'sd35774;
    data[14754] = -'sd77264;
    data[14755] = -'sd49325;
    data[14756] = -'sd17593;
    data[14757] =  'sd40690;
    data[14758] = -'sd42852;
    data[14759] =  'sd27718;
    data[14760] =  'sd30185;
    data[14761] =  'sd47454;
    data[14762] =  'sd4496;
    data[14763] =  'sd31472;
    data[14764] =  'sd56463;
    data[14765] =  'sd67559;
    data[14766] = -'sd18610;
    data[14767] =  'sd33571;
    data[14768] =  'sd71156;
    data[14769] =  'sd6569;
    data[14770] =  'sd45983;
    data[14771] = -'sd5801;
    data[14772] = -'sd40607;
    data[14773] =  'sd43433;
    data[14774] = -'sd23651;
    data[14775] = -'sd1716;
    data[14776] = -'sd12012;
    data[14777] =  'sd79757;
    data[14778] =  'sd66776;
    data[14779] = -'sd24091;
    data[14780] = -'sd4796;
    data[14781] = -'sd33572;
    data[14782] = -'sd71163;
    data[14783] = -'sd6618;
    data[14784] = -'sd46326;
    data[14785] =  'sd3400;
    data[14786] =  'sd23800;
    data[14787] =  'sd2759;
    data[14788] =  'sd19313;
    data[14789] = -'sd28650;
    data[14790] = -'sd36709;
    data[14791] =  'sd70719;
    data[14792] =  'sd3510;
    data[14793] =  'sd24570;
    data[14794] =  'sd8149;
    data[14795] =  'sd57043;
    data[14796] =  'sd71619;
    data[14797] =  'sd9810;
    data[14798] =  'sd68670;
    data[14799] = -'sd10833;
    data[14800] = -'sd75831;
    data[14801] = -'sd39294;
    data[14802] =  'sd52624;
    data[14803] =  'sd40686;
    data[14804] = -'sd42880;
    data[14805] =  'sd27522;
    data[14806] =  'sd28813;
    data[14807] =  'sd37850;
    data[14808] = -'sd62732;
    data[14809] =  'sd52399;
    data[14810] =  'sd39111;
    data[14811] = -'sd53905;
    data[14812] = -'sd49653;
    data[14813] = -'sd19889;
    data[14814] =  'sd24618;
    data[14815] =  'sd8485;
    data[14816] =  'sd59395;
    data[14817] = -'sd75758;
    data[14818] = -'sd38783;
    data[14819] =  'sd56201;
    data[14820] =  'sd65725;
    data[14821] = -'sd31448;
    data[14822] = -'sd56295;
    data[14823] = -'sd66383;
    data[14824] =  'sd26842;
    data[14825] =  'sd24053;
    data[14826] =  'sd4530;
    data[14827] =  'sd31710;
    data[14828] =  'sd58129;
    data[14829] =  'sd79221;
    data[14830] =  'sd63024;
    data[14831] = -'sd50355;
    data[14832] = -'sd24803;
    data[14833] = -'sd9780;
    data[14834] = -'sd68460;
    data[14835] =  'sd12303;
    data[14836] = -'sd77720;
    data[14837] = -'sd52517;
    data[14838] = -'sd39937;
    data[14839] =  'sd48123;
    data[14840] =  'sd9179;
    data[14841] =  'sd64253;
    data[14842] = -'sd41752;
    data[14843] =  'sd35418;
    data[14844] = -'sd79756;
    data[14845] = -'sd66769;
    data[14846] =  'sd24140;
    data[14847] =  'sd5139;
    data[14848] =  'sd35973;
    data[14849] = -'sd75871;
    data[14850] = -'sd39574;
    data[14851] =  'sd50664;
    data[14852] =  'sd26966;
    data[14853] =  'sd24921;
    data[14854] =  'sd10606;
    data[14855] =  'sd74242;
    data[14856] =  'sd28171;
    data[14857] =  'sd33356;
    data[14858] =  'sd69651;
    data[14859] = -'sd3966;
    data[14860] = -'sd27762;
    data[14861] = -'sd30493;
    data[14862] = -'sd49610;
    data[14863] = -'sd19588;
    data[14864] =  'sd26725;
    data[14865] =  'sd23234;
    data[14866] = -'sd1203;
    data[14867] = -'sd8421;
    data[14868] = -'sd58947;
    data[14869] =  'sd78894;
    data[14870] =  'sd60735;
    data[14871] = -'sd66378;
    data[14872] =  'sd26877;
    data[14873] =  'sd24298;
    data[14874] =  'sd6245;
    data[14875] =  'sd43715;
    data[14876] = -'sd21677;
    data[14877] =  'sd12102;
    data[14878] = -'sd79127;
    data[14879] = -'sd62366;
    data[14880] =  'sd54961;
    data[14881] =  'sd57045;
    data[14882] =  'sd71633;
    data[14883] =  'sd9908;
    data[14884] =  'sd69356;
    data[14885] = -'sd6031;
    data[14886] = -'sd42217;
    data[14887] =  'sd32163;
    data[14888] =  'sd61300;
    data[14889] = -'sd62423;
    data[14890] =  'sd54562;
    data[14891] =  'sd54252;
    data[14892] =  'sd52082;
    data[14893] =  'sd36892;
    data[14894] = -'sd69438;
    data[14895] =  'sd5457;
    data[14896] =  'sd38199;
    data[14897] = -'sd60289;
    data[14898] =  'sd69500;
    data[14899] = -'sd5023;
    data[14900] = -'sd35161;
    data[14901] =  'sd81555;
    data[14902] =  'sd79362;
    data[14903] =  'sd64011;
    data[14904] = -'sd43446;
    data[14905] =  'sd23560;
    data[14906] =  'sd1079;
    data[14907] =  'sd7553;
    data[14908] =  'sd52871;
    data[14909] =  'sd42415;
    data[14910] = -'sd30777;
    data[14911] = -'sd51598;
    data[14912] = -'sd33504;
    data[14913] = -'sd70687;
    data[14914] = -'sd3286;
    data[14915] = -'sd23002;
    data[14916] =  'sd2827;
    data[14917] =  'sd19789;
    data[14918] = -'sd25318;
    data[14919] = -'sd13385;
    data[14920] =  'sd70146;
    data[14921] = -'sd501;
    data[14922] = -'sd3507;
    data[14923] = -'sd24549;
    data[14924] = -'sd8002;
    data[14925] = -'sd56014;
    data[14926] = -'sd64416;
    data[14927] =  'sd40611;
    data[14928] = -'sd43405;
    data[14929] =  'sd23847;
    data[14930] =  'sd3088;
    data[14931] =  'sd21616;
    data[14932] = -'sd12529;
    data[14933] =  'sd76138;
    data[14934] =  'sd41443;
    data[14935] = -'sd37581;
    data[14936] =  'sd64615;
    data[14937] = -'sd39218;
    data[14938] =  'sd53156;
    data[14939] =  'sd44410;
    data[14940] = -'sd16812;
    data[14941] =  'sd46157;
    data[14942] = -'sd4583;
    data[14943] = -'sd32081;
    data[14944] = -'sd60726;
    data[14945] =  'sd66441;
    data[14946] = -'sd26436;
    data[14947] = -'sd21211;
    data[14948] =  'sd15364;
    data[14949] = -'sd56293;
    data[14950] = -'sd66369;
    data[14951] =  'sd26940;
    data[14952] =  'sd24739;
    data[14953] =  'sd9332;
    data[14954] =  'sd65324;
    data[14955] = -'sd34255;
    data[14956] = -'sd75944;
    data[14957] = -'sd40085;
    data[14958] =  'sd47087;
    data[14959] =  'sd1927;
    data[14960] =  'sd13489;
    data[14961] = -'sd69418;
    data[14962] =  'sd5597;
    data[14963] =  'sd39179;
    data[14964] = -'sd53429;
    data[14965] = -'sd46321;
    data[14966] =  'sd3435;
    data[14967] =  'sd24045;
    data[14968] =  'sd4474;
    data[14969] =  'sd31318;
    data[14970] =  'sd55385;
    data[14971] =  'sd60013;
    data[14972] = -'sd71432;
    data[14973] = -'sd8501;
    data[14974] = -'sd59507;
    data[14975] =  'sd74974;
    data[14976] =  'sd33295;
    data[14977] =  'sd69224;
    data[14978] = -'sd6955;
    data[14979] = -'sd48685;
    data[14980] = -'sd13113;
    data[14981] =  'sd72050;
    data[14982] =  'sd12827;
    data[14983] = -'sd74052;
    data[14984] = -'sd26841;
    data[14985] = -'sd24046;
    data[14986] = -'sd4481;
    data[14987] = -'sd31367;
    data[14988] = -'sd55728;
    data[14989] = -'sd62414;
    data[14990] =  'sd54625;
    data[14991] =  'sd54693;
    data[14992] =  'sd55169;
    data[14993] =  'sd58501;
    data[14994] =  'sd81825;
    data[14995] =  'sd81252;
    data[14996] =  'sd77241;
    data[14997] =  'sd49164;
    data[14998] =  'sd16466;
    data[14999] = -'sd48579;
    data[15000] = -'sd12371;
    data[15001] =  'sd77244;
    data[15002] =  'sd49185;
    data[15003] =  'sd16613;
    data[15004] = -'sd47550;
    data[15005] = -'sd5168;
    data[15006] = -'sd36176;
    data[15007] =  'sd74450;
    data[15008] =  'sd29627;
    data[15009] =  'sd43548;
    data[15010] = -'sd22846;
    data[15011] =  'sd3919;
    data[15012] =  'sd27433;
    data[15013] =  'sd28190;
    data[15014] =  'sd33489;
    data[15015] =  'sd70582;
    data[15016] =  'sd2551;
    data[15017] =  'sd17857;
    data[15018] = -'sd38842;
    data[15019] =  'sd55788;
    data[15020] =  'sd62834;
    data[15021] = -'sd51685;
    data[15022] = -'sd34113;
    data[15023] = -'sd74950;
    data[15024] = -'sd33127;
    data[15025] = -'sd68048;
    data[15026] =  'sd15187;
    data[15027] = -'sd57532;
    data[15028] = -'sd75042;
    data[15029] = -'sd33771;
    data[15030] = -'sd72556;
    data[15031] = -'sd16369;
    data[15032] =  'sd49258;
    data[15033] =  'sd17124;
    data[15034] = -'sd43973;
    data[15035] =  'sd19871;
    data[15036] = -'sd24744;
    data[15037] = -'sd9367;
    data[15038] = -'sd65569;
    data[15039] =  'sd32540;
    data[15040] =  'sd63939;
    data[15041] = -'sd43950;
    data[15042] =  'sd20032;
    data[15043] = -'sd23617;
    data[15044] = -'sd1478;
    data[15045] = -'sd10346;
    data[15046] = -'sd72422;
    data[15047] = -'sd15431;
    data[15048] =  'sd55824;
    data[15049] =  'sd63086;
    data[15050] = -'sd49921;
    data[15051] = -'sd21765;
    data[15052] =  'sd11486;
    data[15053] =  'sd80402;
    data[15054] =  'sd71291;
    data[15055] =  'sd7514;
    data[15056] =  'sd52598;
    data[15057] =  'sd40504;
    data[15058] = -'sd44154;
    data[15059] =  'sd18604;
    data[15060] = -'sd33613;
    data[15061] = -'sd71450;
    data[15062] = -'sd8627;
    data[15063] = -'sd60389;
    data[15064] =  'sd68800;
    data[15065] = -'sd9923;
    data[15066] = -'sd69461;
    data[15067] =  'sd5296;
    data[15068] =  'sd37072;
    data[15069] = -'sd68178;
    data[15070] =  'sd14277;
    data[15071] = -'sd63902;
    data[15072] =  'sd44209;
    data[15073] = -'sd18219;
    data[15074] =  'sd36308;
    data[15075] = -'sd73526;
    data[15076] = -'sd23159;
    data[15077] =  'sd1728;
    data[15078] =  'sd12096;
    data[15079] = -'sd79169;
    data[15080] = -'sd62660;
    data[15081] =  'sd52903;
    data[15082] =  'sd42639;
    data[15083] = -'sd29209;
    data[15084] = -'sd40622;
    data[15085] =  'sd43328;
    data[15086] = -'sd24386;
    data[15087] = -'sd6861;
    data[15088] = -'sd48027;
    data[15089] = -'sd8507;
    data[15090] = -'sd59549;
    data[15091] =  'sd74680;
    data[15092] =  'sd31237;
    data[15093] =  'sd54818;
    data[15094] =  'sd56044;
    data[15095] =  'sd64626;
    data[15096] = -'sd39141;
    data[15097] =  'sd53695;
    data[15098] =  'sd48183;
    data[15099] =  'sd9599;
    data[15100] =  'sd67193;
    data[15101] = -'sd21172;
    data[15102] =  'sd15637;
    data[15103] = -'sd54382;
    data[15104] = -'sd52992;
    data[15105] = -'sd43262;
    data[15106] =  'sd24848;
    data[15107] =  'sd10095;
    data[15108] =  'sd70665;
    data[15109] =  'sd3132;
    data[15110] =  'sd21924;
    data[15111] = -'sd10373;
    data[15112] = -'sd72611;
    data[15113] = -'sd16754;
    data[15114] =  'sd46563;
    data[15115] = -'sd1741;
    data[15116] = -'sd12187;
    data[15117] =  'sd78532;
    data[15118] =  'sd58201;
    data[15119] =  'sd79725;
    data[15120] =  'sd66552;
    data[15121] = -'sd25659;
    data[15122] = -'sd15772;
    data[15123] =  'sd53437;
    data[15124] =  'sd46377;
    data[15125] = -'sd3043;
    data[15126] = -'sd21301;
    data[15127] =  'sd14734;
    data[15128] = -'sd60703;
    data[15129] =  'sd66602;
    data[15130] = -'sd25309;
    data[15131] = -'sd13322;
    data[15132] =  'sd70587;
    data[15133] =  'sd2586;
    data[15134] =  'sd18102;
    data[15135] = -'sd37127;
    data[15136] =  'sd67793;
    data[15137] = -'sd16972;
    data[15138] =  'sd45037;
    data[15139] = -'sd12423;
    data[15140] =  'sd76880;
    data[15141] =  'sd46637;
    data[15142] = -'sd1223;
    data[15143] = -'sd8561;
    data[15144] = -'sd59927;
    data[15145] =  'sd72034;
    data[15146] =  'sd12715;
    data[15147] = -'sd74836;
    data[15148] = -'sd32329;
    data[15149] = -'sd62462;
    data[15150] =  'sd54289;
    data[15151] =  'sd52341;
    data[15152] =  'sd38705;
    data[15153] = -'sd56747;
    data[15154] = -'sd69547;
    data[15155] =  'sd4694;
    data[15156] =  'sd32858;
    data[15157] =  'sd66165;
    data[15158] = -'sd28368;
    data[15159] = -'sd34735;
    data[15160] = -'sd79304;
    data[15161] = -'sd63605;
    data[15162] =  'sd46288;
    data[15163] = -'sd3666;
    data[15164] = -'sd25662;
    data[15165] = -'sd15793;
    data[15166] =  'sd53290;
    data[15167] =  'sd45348;
    data[15168] = -'sd10246;
    data[15169] = -'sd71722;
    data[15170] = -'sd10531;
    data[15171] = -'sd73717;
    data[15172] = -'sd24496;
    data[15173] = -'sd7631;
    data[15174] = -'sd53417;
    data[15175] = -'sd46237;
    data[15176] =  'sd4023;
    data[15177] =  'sd28161;
    data[15178] =  'sd33286;
    data[15179] =  'sd69161;
    data[15180] = -'sd7396;
    data[15181] = -'sd51772;
    data[15182] = -'sd34722;
    data[15183] = -'sd79213;
    data[15184] = -'sd62968;
    data[15185] =  'sd50747;
    data[15186] =  'sd27547;
    data[15187] =  'sd28988;
    data[15188] =  'sd39075;
    data[15189] = -'sd54157;
    data[15190] = -'sd51417;
    data[15191] = -'sd32237;
    data[15192] = -'sd61818;
    data[15193] =  'sd58797;
    data[15194] = -'sd79944;
    data[15195] = -'sd68085;
    data[15196] =  'sd14928;
    data[15197] = -'sd59345;
    data[15198] =  'sd76108;
    data[15199] =  'sd41233;
    data[15200] = -'sd39051;
    data[15201] =  'sd54325;
    data[15202] =  'sd52593;
    data[15203] =  'sd40469;
    data[15204] = -'sd44399;
    data[15205] =  'sd16889;
    data[15206] = -'sd45618;
    data[15207] =  'sd8356;
    data[15208] =  'sd58492;
    data[15209] =  'sd81762;
    data[15210] =  'sd80811;
    data[15211] =  'sd74154;
    data[15212] =  'sd27555;
    data[15213] =  'sd29044;
    data[15214] =  'sd39467;
    data[15215] = -'sd51413;
    data[15216] = -'sd32209;
    data[15217] = -'sd61622;
    data[15218] =  'sd60169;
    data[15219] = -'sd70340;
    data[15220] = -'sd857;
    data[15221] = -'sd5999;
    data[15222] = -'sd41993;
    data[15223] =  'sd33731;
    data[15224] =  'sd72276;
    data[15225] =  'sd14409;
    data[15226] = -'sd62978;
    data[15227] =  'sd50677;
    data[15228] =  'sd27057;
    data[15229] =  'sd25558;
    data[15230] =  'sd15065;
    data[15231] = -'sd58386;
    data[15232] = -'sd81020;
    data[15233] = -'sd75617;
    data[15234] = -'sd37796;
    data[15235] =  'sd63110;
    data[15236] = -'sd49753;
    data[15237] = -'sd20589;
    data[15238] =  'sd19718;
    data[15239] = -'sd25815;
    data[15240] = -'sd16864;
    data[15241] =  'sd45793;
    data[15242] = -'sd7131;
    data[15243] = -'sd49917;
    data[15244] = -'sd21737;
    data[15245] =  'sd11682;
    data[15246] =  'sd81774;
    data[15247] =  'sd80895;
    data[15248] =  'sd74742;
    data[15249] =  'sd31671;
    data[15250] =  'sd57856;
    data[15251] =  'sd77310;
    data[15252] =  'sd49647;
    data[15253] =  'sd19847;
    data[15254] = -'sd24912;
    data[15255] = -'sd10543;
    data[15256] = -'sd73801;
    data[15257] = -'sd25084;
    data[15258] = -'sd11747;
    data[15259] =  'sd81612;
    data[15260] =  'sd79761;
    data[15261] =  'sd66804;
    data[15262] = -'sd23895;
    data[15263] = -'sd3424;
    data[15264] = -'sd23968;
    data[15265] = -'sd3935;
    data[15266] = -'sd27545;
    data[15267] = -'sd28974;
    data[15268] = -'sd38977;
    data[15269] =  'sd54843;
    data[15270] =  'sd56219;
    data[15271] =  'sd65851;
    data[15272] = -'sd30566;
    data[15273] = -'sd50121;
    data[15274] = -'sd23165;
    data[15275] =  'sd1686;
    data[15276] =  'sd11802;
    data[15277] = -'sd81227;
    data[15278] = -'sd77066;
    data[15279] = -'sd47939;
    data[15280] = -'sd7891;
    data[15281] = -'sd55237;
    data[15282] = -'sd58977;
    data[15283] =  'sd78684;
    data[15284] =  'sd59265;
    data[15285] = -'sd76668;
    data[15286] = -'sd45153;
    data[15287] =  'sd11611;
    data[15288] =  'sd81277;
    data[15289] =  'sd77416;
    data[15290] =  'sd50389;
    data[15291] =  'sd25041;
    data[15292] =  'sd11446;
    data[15293] =  'sd80122;
    data[15294] =  'sd69331;
    data[15295] = -'sd6206;
    data[15296] = -'sd43442;
    data[15297] =  'sd23588;
    data[15298] =  'sd1275;
    data[15299] =  'sd8925;
    data[15300] =  'sd62475;
    data[15301] = -'sd54198;
    data[15302] = -'sd51704;
    data[15303] = -'sd34246;
    data[15304] = -'sd75881;
    data[15305] = -'sd39644;
    data[15306] =  'sd50174;
    data[15307] =  'sd23536;
    data[15308] =  'sd911;
    data[15309] =  'sd6377;
    data[15310] =  'sd44639;
    data[15311] = -'sd15209;
    data[15312] =  'sd57378;
    data[15313] =  'sd73964;
    data[15314] =  'sd26225;
    data[15315] =  'sd19734;
    data[15316] = -'sd25703;
    data[15317] = -'sd16080;
    data[15318] =  'sd51281;
    data[15319] =  'sd31285;
    data[15320] =  'sd55154;
    data[15321] =  'sd58396;
    data[15322] =  'sd81090;
    data[15323] =  'sd76107;
    data[15324] =  'sd41226;
    data[15325] = -'sd39100;
    data[15326] =  'sd53982;
    data[15327] =  'sd50192;
    data[15328] =  'sd23662;
    data[15329] =  'sd1793;
    data[15330] =  'sd12551;
    data[15331] = -'sd75984;
    data[15332] = -'sd40365;
    data[15333] =  'sd45127;
    data[15334] = -'sd11793;
    data[15335] =  'sd81290;
    data[15336] =  'sd77507;
    data[15337] =  'sd51026;
    data[15338] =  'sd29500;
    data[15339] =  'sd42659;
    data[15340] = -'sd29069;
    data[15341] = -'sd39642;
    data[15342] =  'sd50188;
    data[15343] =  'sd23634;
    data[15344] =  'sd1597;
    data[15345] =  'sd11179;
    data[15346] =  'sd78253;
    data[15347] =  'sd56248;
    data[15348] =  'sd66054;
    data[15349] = -'sd29145;
    data[15350] = -'sd40174;
    data[15351] =  'sd46464;
    data[15352] = -'sd2434;
    data[15353] = -'sd17038;
    data[15354] =  'sd44575;
    data[15355] = -'sd15657;
    data[15356] =  'sd54242;
    data[15357] =  'sd52012;
    data[15358] =  'sd36402;
    data[15359] = -'sd72868;
    data[15360] = -'sd18553;
    data[15361] =  'sd33970;
    data[15362] =  'sd73949;
    data[15363] =  'sd26120;
    data[15364] =  'sd18999;
    data[15365] = -'sd30848;
    data[15366] = -'sd52095;
    data[15367] = -'sd36983;
    data[15368] =  'sd68801;
    data[15369] = -'sd9916;
    data[15370] = -'sd69412;
    data[15371] =  'sd5639;
    data[15372] =  'sd39473;
    data[15373] = -'sd51371;
    data[15374] = -'sd31915;
    data[15375] = -'sd59564;
    data[15376] =  'sd74575;
    data[15377] =  'sd30502;
    data[15378] =  'sd49673;
    data[15379] =  'sd20029;
    data[15380] = -'sd23638;
    data[15381] = -'sd1625;
    data[15382] = -'sd11375;
    data[15383] = -'sd79625;
    data[15384] = -'sd65852;
    data[15385] =  'sd30559;
    data[15386] =  'sd50072;
    data[15387] =  'sd22822;
    data[15388] = -'sd4087;
    data[15389] = -'sd28609;
    data[15390] = -'sd36422;
    data[15391] =  'sd72728;
    data[15392] =  'sd17573;
    data[15393] = -'sd40830;
    data[15394] =  'sd41872;
    data[15395] = -'sd34578;
    data[15396] = -'sd78205;
    data[15397] = -'sd55912;
    data[15398] = -'sd63702;
    data[15399] =  'sd45609;
    data[15400] = -'sd8419;
    data[15401] = -'sd58933;
    data[15402] =  'sd78992;
    data[15403] =  'sd61421;
    data[15404] = -'sd61576;
    data[15405] =  'sd60491;
    data[15406] = -'sd68086;
    data[15407] =  'sd14921;
    data[15408] = -'sd59394;
    data[15409] =  'sd75765;
    data[15410] =  'sd38832;
    data[15411] = -'sd55858;
    data[15412] = -'sd63324;
    data[15413] =  'sd48255;
    data[15414] =  'sd10103;
    data[15415] =  'sd70721;
    data[15416] =  'sd3524;
    data[15417] =  'sd24668;
    data[15418] =  'sd8835;
    data[15419] =  'sd61845;
    data[15420] = -'sd58608;
    data[15421] =  'sd81267;
    data[15422] =  'sd77346;
    data[15423] =  'sd49899;
    data[15424] =  'sd21611;
    data[15425] = -'sd12564;
    data[15426] =  'sd75893;
    data[15427] =  'sd39728;
    data[15428] = -'sd49586;
    data[15429] = -'sd19420;
    data[15430] =  'sd27901;
    data[15431] =  'sd31466;
    data[15432] =  'sd56421;
    data[15433] =  'sd67265;
    data[15434] = -'sd20668;
    data[15435] =  'sd19165;
    data[15436] = -'sd29686;
    data[15437] = -'sd43961;
    data[15438] =  'sd19955;
    data[15439] = -'sd24156;
    data[15440] = -'sd5251;
    data[15441] = -'sd36757;
    data[15442] =  'sd70383;
    data[15443] =  'sd1158;
    data[15444] =  'sd8106;
    data[15445] =  'sd56742;
    data[15446] =  'sd69512;
    data[15447] = -'sd4939;
    data[15448] = -'sd34573;
    data[15449] = -'sd78170;
    data[15450] = -'sd55667;
    data[15451] = -'sd61987;
    data[15452] =  'sd57614;
    data[15453] =  'sd75616;
    data[15454] =  'sd37789;
    data[15455] = -'sd63159;
    data[15456] =  'sd49410;
    data[15457] =  'sd18188;
    data[15458] = -'sd36525;
    data[15459] =  'sd72007;
    data[15460] =  'sd12526;
    data[15461] = -'sd76159;
    data[15462] = -'sd41590;
    data[15463] =  'sd36552;
    data[15464] = -'sd71818;
    data[15465] = -'sd11203;
    data[15466] = -'sd78421;
    data[15467] = -'sd57424;
    data[15468] = -'sd74286;
    data[15469] = -'sd28479;
    data[15470] = -'sd35512;
    data[15471] =  'sd79098;
    data[15472] =  'sd62163;
    data[15473] = -'sd56382;
    data[15474] = -'sd66992;
    data[15475] =  'sd22579;
    data[15476] = -'sd5788;
    data[15477] = -'sd40516;
    data[15478] =  'sd44070;
    data[15479] = -'sd19192;
    data[15480] =  'sd29497;
    data[15481] =  'sd42638;
    data[15482] = -'sd29216;
    data[15483] = -'sd40671;
    data[15484] =  'sd42985;
    data[15485] = -'sd26787;
    data[15486] = -'sd23668;
    data[15487] = -'sd1835;
    data[15488] = -'sd12845;
    data[15489] =  'sd73926;
    data[15490] =  'sd25959;
    data[15491] =  'sd17872;
    data[15492] = -'sd38737;
    data[15493] =  'sd56523;
    data[15494] =  'sd67979;
    data[15495] = -'sd15670;
    data[15496] =  'sd54151;
    data[15497] =  'sd51375;
    data[15498] =  'sd31943;
    data[15499] =  'sd59760;
    data[15500] = -'sd73203;
    data[15501] = -'sd20898;
    data[15502] =  'sd17555;
    data[15503] = -'sd40956;
    data[15504] =  'sd40990;
    data[15505] = -'sd40752;
    data[15506] =  'sd42418;
    data[15507] = -'sd30756;
    data[15508] = -'sd51451;
    data[15509] = -'sd32475;
    data[15510] = -'sd63484;
    data[15511] =  'sd47135;
    data[15512] =  'sd2263;
    data[15513] =  'sd15841;
    data[15514] = -'sd52954;
    data[15515] = -'sd42996;
    data[15516] =  'sd26710;
    data[15517] =  'sd23129;
    data[15518] = -'sd1938;
    data[15519] = -'sd13566;
    data[15520] =  'sd68879;
    data[15521] = -'sd9370;
    data[15522] = -'sd65590;
    data[15523] =  'sd32393;
    data[15524] =  'sd62910;
    data[15525] = -'sd51153;
    data[15526] = -'sd30389;
    data[15527] = -'sd48882;
    data[15528] = -'sd14492;
    data[15529] =  'sd62397;
    data[15530] = -'sd54744;
    data[15531] = -'sd55526;
    data[15532] = -'sd61000;
    data[15533] =  'sd64523;
    data[15534] = -'sd39862;
    data[15535] =  'sd48648;
    data[15536] =  'sd12854;
    data[15537] = -'sd73863;
    data[15538] = -'sd25518;
    data[15539] = -'sd14785;
    data[15540] =  'sd60346;
    data[15541] = -'sd69101;
    data[15542] =  'sd7816;
    data[15543] =  'sd54712;
    data[15544] =  'sd55302;
    data[15545] =  'sd59432;
    data[15546] = -'sd75499;
    data[15547] = -'sd36970;
    data[15548] =  'sd68892;
    data[15549] = -'sd9279;
    data[15550] = -'sd64953;
    data[15551] =  'sd36852;
    data[15552] = -'sd69718;
    data[15553] =  'sd3497;
    data[15554] =  'sd24479;
    data[15555] =  'sd7512;
    data[15556] =  'sd52584;
    data[15557] =  'sd40406;
    data[15558] = -'sd44840;
    data[15559] =  'sd13802;
    data[15560] = -'sd67227;
    data[15561] =  'sd20934;
    data[15562] = -'sd17303;
    data[15563] =  'sd42720;
    data[15564] = -'sd28642;
    data[15565] = -'sd36653;
    data[15566] =  'sd71111;
    data[15567] =  'sd6254;
    data[15568] =  'sd43778;
    data[15569] = -'sd21236;
    data[15570] =  'sd15189;
    data[15571] = -'sd57518;
    data[15572] = -'sd74944;
    data[15573] = -'sd33085;
    data[15574] = -'sd67754;
    data[15575] =  'sd17245;
    data[15576] = -'sd43126;
    data[15577] =  'sd25800;
    data[15578] =  'sd16759;
    data[15579] = -'sd46528;
    data[15580] =  'sd1986;
    data[15581] =  'sd13902;
    data[15582] = -'sd66527;
    data[15583] =  'sd25834;
    data[15584] =  'sd16997;
    data[15585] = -'sd44862;
    data[15586] =  'sd13648;
    data[15587] = -'sd68305;
    data[15588] =  'sd13388;
    data[15589] = -'sd70125;
    data[15590] =  'sd648;
    data[15591] =  'sd4536;
    data[15592] =  'sd31752;
    data[15593] =  'sd58423;
    data[15594] =  'sd81279;
    data[15595] =  'sd77430;
    data[15596] =  'sd50487;
    data[15597] =  'sd25727;
    data[15598] =  'sd16248;
    data[15599] = -'sd50105;
    data[15600] = -'sd23053;
    data[15601] =  'sd2470;
    data[15602] =  'sd17290;
    data[15603] = -'sd42811;
    data[15604] =  'sd28005;
    data[15605] =  'sd32194;
    data[15606] =  'sd61517;
    data[15607] = -'sd60904;
    data[15608] =  'sd65195;
    data[15609] = -'sd35158;
    data[15610] =  'sd81576;
    data[15611] =  'sd79509;
    data[15612] =  'sd65040;
    data[15613] = -'sd36243;
    data[15614] =  'sd73981;
    data[15615] =  'sd26344;
    data[15616] =  'sd20567;
    data[15617] = -'sd19872;
    data[15618] =  'sd24737;
    data[15619] =  'sd9318;
    data[15620] =  'sd65226;
    data[15621] = -'sd34941;
    data[15622] = -'sd80746;
    data[15623] = -'sd73699;
    data[15624] = -'sd24370;
    data[15625] = -'sd6749;
    data[15626] = -'sd47243;
    data[15627] = -'sd3019;
    data[15628] = -'sd21133;
    data[15629] =  'sd15910;
    data[15630] = -'sd52471;
    data[15631] = -'sd39615;
    data[15632] =  'sd50377;
    data[15633] =  'sd24957;
    data[15634] =  'sd10858;
    data[15635] =  'sd76006;
    data[15636] =  'sd40519;
    data[15637] = -'sd44049;
    data[15638] =  'sd19339;
    data[15639] = -'sd28468;
    data[15640] = -'sd35435;
    data[15641] =  'sd79637;
    data[15642] =  'sd65936;
    data[15643] = -'sd29971;
    data[15644] = -'sd45956;
    data[15645] =  'sd5990;
    data[15646] =  'sd41930;
    data[15647] = -'sd34172;
    data[15648] = -'sd75363;
    data[15649] = -'sd36018;
    data[15650] =  'sd75556;
    data[15651] =  'sd37369;
    data[15652] = -'sd66099;
    data[15653] =  'sd28830;
    data[15654] =  'sd37969;
    data[15655] = -'sd61899;
    data[15656] =  'sd58230;
    data[15657] =  'sd79928;
    data[15658] =  'sd67973;
    data[15659] = -'sd15712;
    data[15660] =  'sd53857;
    data[15661] =  'sd49317;
    data[15662] =  'sd17537;
    data[15663] = -'sd41082;
    data[15664] =  'sd40108;
    data[15665] = -'sd46926;
    data[15666] = -'sd800;
    data[15667] = -'sd5600;
    data[15668] = -'sd39200;
    data[15669] =  'sd53282;
    data[15670] =  'sd45292;
    data[15671] = -'sd10638;
    data[15672] = -'sd74466;
    data[15673] = -'sd29739;
    data[15674] = -'sd44332;
    data[15675] =  'sd17358;
    data[15676] = -'sd42335;
    data[15677] =  'sd31337;
    data[15678] =  'sd55518;
    data[15679] =  'sd60944;
    data[15680] = -'sd64915;
    data[15681] =  'sd37118;
    data[15682] = -'sd67856;
    data[15683] =  'sd16531;
    data[15684] = -'sd48124;
    data[15685] = -'sd9186;
    data[15686] = -'sd64302;
    data[15687] =  'sd41409;
    data[15688] = -'sd37819;
    data[15689] =  'sd62949;
    data[15690] = -'sd50880;
    data[15691] = -'sd28478;
    data[15692] = -'sd35505;
    data[15693] =  'sd79147;
    data[15694] =  'sd62506;
    data[15695] = -'sd53981;
    data[15696] = -'sd50185;
    data[15697] = -'sd23613;
    data[15698] = -'sd1450;
    data[15699] = -'sd10150;
    data[15700] = -'sd71050;
    data[15701] = -'sd5827;
    data[15702] = -'sd40789;
    data[15703] =  'sd42159;
    data[15704] = -'sd32569;
    data[15705] = -'sd64142;
    data[15706] =  'sd42529;
    data[15707] = -'sd29979;
    data[15708] = -'sd46012;
    data[15709] =  'sd5598;
    data[15710] =  'sd39186;
    data[15711] = -'sd53380;
    data[15712] = -'sd45978;
    data[15713] =  'sd5836;
    data[15714] =  'sd40852;
    data[15715] = -'sd41718;
    data[15716] =  'sd35656;
    data[15717] = -'sd78090;
    data[15718] = -'sd55107;
    data[15719] = -'sd58067;
    data[15720] = -'sd78787;
    data[15721] = -'sd59986;
    data[15722] =  'sd71621;
    data[15723] =  'sd9824;
    data[15724] =  'sd68768;
    data[15725] = -'sd10147;
    data[15726] = -'sd71029;
    data[15727] = -'sd5680;
    data[15728] = -'sd39760;
    data[15729] =  'sd49362;
    data[15730] =  'sd17852;
    data[15731] = -'sd38877;
    data[15732] =  'sd55543;
    data[15733] =  'sd61119;
    data[15734] = -'sd63690;
    data[15735] =  'sd45693;
    data[15736] = -'sd7831;
    data[15737] = -'sd54817;
    data[15738] = -'sd56037;
    data[15739] = -'sd64577;
    data[15740] =  'sd39484;
    data[15741] = -'sd51294;
    data[15742] = -'sd31376;
    data[15743] = -'sd55791;
    data[15744] = -'sd62855;
    data[15745] =  'sd51538;
    data[15746] =  'sd33084;
    data[15747] =  'sd67747;
    data[15748] = -'sd17294;
    data[15749] =  'sd42783;
    data[15750] = -'sd28201;
    data[15751] = -'sd33566;
    data[15752] = -'sd71121;
    data[15753] = -'sd6324;
    data[15754] = -'sd44268;
    data[15755] =  'sd17806;
    data[15756] = -'sd39199;
    data[15757] =  'sd53289;
    data[15758] =  'sd45341;
    data[15759] = -'sd10295;
    data[15760] = -'sd72065;
    data[15761] = -'sd12932;
    data[15762] =  'sd73317;
    data[15763] =  'sd21696;
    data[15764] = -'sd11969;
    data[15765] =  'sd80058;
    data[15766] =  'sd68883;
    data[15767] = -'sd9342;
    data[15768] = -'sd65394;
    data[15769] =  'sd33765;
    data[15770] =  'sd72514;
    data[15771] =  'sd16075;
    data[15772] = -'sd51316;
    data[15773] = -'sd31530;
    data[15774] = -'sd56869;
    data[15775] = -'sd70401;
    data[15776] = -'sd1284;
    data[15777] = -'sd8988;
    data[15778] = -'sd62916;
    data[15779] =  'sd51111;
    data[15780] =  'sd30095;
    data[15781] =  'sd46824;
    data[15782] =  'sd86;
    data[15783] =  'sd602;
    data[15784] =  'sd4214;
    data[15785] =  'sd29498;
    data[15786] =  'sd42645;
    data[15787] = -'sd29167;
    data[15788] = -'sd40328;
    data[15789] =  'sd45386;
    data[15790] = -'sd9980;
    data[15791] = -'sd69860;
    data[15792] =  'sd2503;
    data[15793] =  'sd17521;
    data[15794] = -'sd41194;
    data[15795] =  'sd39324;
    data[15796] = -'sd52414;
    data[15797] = -'sd39216;
    data[15798] =  'sd53170;
    data[15799] =  'sd44508;
    data[15800] = -'sd16126;
    data[15801] =  'sd50959;
    data[15802] =  'sd29031;
    data[15803] =  'sd39376;
    data[15804] = -'sd52050;
    data[15805] = -'sd36668;
    data[15806] =  'sd71006;
    data[15807] =  'sd5519;
    data[15808] =  'sd38633;
    data[15809] = -'sd57251;
    data[15810] = -'sd73075;
    data[15811] = -'sd20002;
    data[15812] =  'sd23827;
    data[15813] =  'sd2948;
    data[15814] =  'sd20636;
    data[15815] = -'sd19389;
    data[15816] =  'sd28118;
    data[15817] =  'sd32985;
    data[15818] =  'sd67054;
    data[15819] = -'sd22145;
    data[15820] =  'sd8826;
    data[15821] =  'sd61782;
    data[15822] = -'sd59049;
    data[15823] =  'sd78180;
    data[15824] =  'sd55737;
    data[15825] =  'sd62477;
    data[15826] = -'sd54184;
    data[15827] = -'sd51606;
    data[15828] = -'sd33560;
    data[15829] = -'sd71079;
    data[15830] = -'sd6030;
    data[15831] = -'sd42210;
    data[15832] =  'sd32212;
    data[15833] =  'sd61643;
    data[15834] = -'sd60022;
    data[15835] =  'sd71369;
    data[15836] =  'sd8060;
    data[15837] =  'sd56420;
    data[15838] =  'sd67258;
    data[15839] = -'sd20717;
    data[15840] =  'sd18822;
    data[15841] = -'sd32087;
    data[15842] = -'sd60768;
    data[15843] =  'sd66147;
    data[15844] = -'sd28494;
    data[15845] = -'sd35617;
    data[15846] =  'sd78363;
    data[15847] =  'sd57018;
    data[15848] =  'sd71444;
    data[15849] =  'sd8585;
    data[15850] =  'sd60095;
    data[15851] = -'sd70858;
    data[15852] = -'sd4483;
    data[15853] = -'sd31381;
    data[15854] = -'sd55826;
    data[15855] = -'sd63100;
    data[15856] =  'sd49823;
    data[15857] =  'sd21079;
    data[15858] = -'sd16288;
    data[15859] =  'sd49825;
    data[15860] =  'sd21093;
    data[15861] = -'sd16190;
    data[15862] =  'sd50511;
    data[15863] =  'sd25895;
    data[15864] =  'sd17424;
    data[15865] = -'sd41873;
    data[15866] =  'sd34571;
    data[15867] =  'sd78156;
    data[15868] =  'sd55569;
    data[15869] =  'sd61301;
    data[15870] = -'sd62416;
    data[15871] =  'sd54611;
    data[15872] =  'sd54595;
    data[15873] =  'sd54483;
    data[15874] =  'sd53699;
    data[15875] =  'sd48211;
    data[15876] =  'sd9795;
    data[15877] =  'sd68565;
    data[15878] = -'sd11568;
    data[15879] = -'sd80976;
    data[15880] = -'sd75309;
    data[15881] = -'sd35640;
    data[15882] =  'sd78202;
    data[15883] =  'sd55891;
    data[15884] =  'sd63555;
    data[15885] = -'sd46638;
    data[15886] =  'sd1216;
    data[15887] =  'sd8512;
    data[15888] =  'sd59584;
    data[15889] = -'sd74435;
    data[15890] = -'sd29522;
    data[15891] = -'sd42813;
    data[15892] =  'sd27991;
    data[15893] =  'sd32096;
    data[15894] =  'sd60831;
    data[15895] = -'sd65706;
    data[15896] =  'sd31581;
    data[15897] =  'sd57226;
    data[15898] =  'sd72900;
    data[15899] =  'sd18777;
    data[15900] = -'sd32402;
    data[15901] = -'sd62973;
    data[15902] =  'sd50712;
    data[15903] =  'sd27302;
    data[15904] =  'sd27273;
    data[15905] =  'sd27070;
    data[15906] =  'sd25649;
    data[15907] =  'sd15702;
    data[15908] = -'sd53927;
    data[15909] = -'sd49807;
    data[15910] = -'sd20967;
    data[15911] =  'sd17072;
    data[15912] = -'sd44337;
    data[15913] =  'sd17323;
    data[15914] = -'sd42580;
    data[15915] =  'sd29622;
    data[15916] =  'sd43513;
    data[15917] = -'sd23091;
    data[15918] =  'sd2204;
    data[15919] =  'sd15428;
    data[15920] = -'sd55845;
    data[15921] = -'sd63233;
    data[15922] =  'sd48892;
    data[15923] =  'sd14562;
    data[15924] = -'sd61907;
    data[15925] =  'sd58174;
    data[15926] =  'sd79536;
    data[15927] =  'sd65229;
    data[15928] = -'sd34920;
    data[15929] = -'sd80599;
    data[15930] = -'sd72670;
    data[15931] = -'sd17167;
    data[15932] =  'sd43672;
    data[15933] = -'sd21978;
    data[15934] =  'sd9995;
    data[15935] =  'sd69965;
    data[15936] = -'sd1768;
    data[15937] = -'sd12376;
    data[15938] =  'sd77209;
    data[15939] =  'sd48940;
    data[15940] =  'sd14898;
    data[15941] = -'sd59555;
    data[15942] =  'sd74638;
    data[15943] =  'sd30943;
    data[15944] =  'sd52760;
    data[15945] =  'sd41638;
    data[15946] = -'sd36216;
    data[15947] =  'sd74170;
    data[15948] =  'sd27667;
    data[15949] =  'sd29828;
    data[15950] =  'sd44955;
    data[15951] = -'sd12997;
    data[15952] =  'sd72862;
    data[15953] =  'sd18511;
    data[15954] = -'sd34264;
    data[15955] = -'sd76007;
    data[15956] = -'sd40526;
    data[15957] =  'sd44000;
    data[15958] = -'sd19682;
    data[15959] =  'sd26067;
    data[15960] =  'sd18628;
    data[15961] = -'sd33445;
    data[15962] = -'sd70274;
    data[15963] = -'sd395;
    data[15964] = -'sd2765;
    data[15965] = -'sd19355;
    data[15966] =  'sd28356;
    data[15967] =  'sd34651;
    data[15968] =  'sd78716;
    data[15969] =  'sd59489;
    data[15970] = -'sd75100;
    data[15971] = -'sd34177;
    data[15972] = -'sd75398;
    data[15973] = -'sd36263;
    data[15974] =  'sd73841;
    data[15975] =  'sd25364;
    data[15976] =  'sd13707;
    data[15977] = -'sd67892;
    data[15978] =  'sd16279;
    data[15979] = -'sd49888;
    data[15980] = -'sd21534;
    data[15981] =  'sd13103;
    data[15982] = -'sd72120;
    data[15983] = -'sd13317;
    data[15984] =  'sd70622;
    data[15985] =  'sd2831;
    data[15986] =  'sd19817;
    data[15987] = -'sd25122;
    data[15988] = -'sd12013;
    data[15989] =  'sd79750;
    data[15990] =  'sd66727;
    data[15991] = -'sd24434;
    data[15992] = -'sd7197;
    data[15993] = -'sd50379;
    data[15994] = -'sd24971;
    data[15995] = -'sd10956;
    data[15996] = -'sd76692;
    data[15997] = -'sd45321;
    data[15998] =  'sd10435;
    data[15999] =  'sd73045;
    data[16000] =  'sd19792;
    data[16001] = -'sd25297;
    data[16002] = -'sd13238;
    data[16003] =  'sd71175;
    data[16004] =  'sd6702;
    data[16005] =  'sd46914;
    data[16006] =  'sd716;
    data[16007] =  'sd5012;
    data[16008] =  'sd35084;
    data[16009] =  'sd81747;
    data[16010] =  'sd80706;
    data[16011] =  'sd73419;
    data[16012] =  'sd22410;
    data[16013] = -'sd6971;
    data[16014] = -'sd48797;
    data[16015] = -'sd13897;
    data[16016] =  'sd66562;
    data[16017] = -'sd25589;
    data[16018] = -'sd15282;
    data[16019] =  'sd56867;
    data[16020] =  'sd70387;
    data[16021] =  'sd1186;
    data[16022] =  'sd8302;
    data[16023] =  'sd58114;
    data[16024] =  'sd79116;
    data[16025] =  'sd62289;
    data[16026] = -'sd55500;
    data[16027] = -'sd60818;
    data[16028] =  'sd65797;
    data[16029] = -'sd30944;
    data[16030] = -'sd52767;
    data[16031] = -'sd41687;
    data[16032] =  'sd35873;
    data[16033] = -'sd76571;
    data[16034] = -'sd44474;
    data[16035] =  'sd16364;
    data[16036] = -'sd49293;
    data[16037] = -'sd17369;
    data[16038] =  'sd42258;
    data[16039] = -'sd31876;
    data[16040] = -'sd59291;
    data[16041] =  'sd76486;
    data[16042] =  'sd43879;
    data[16043] = -'sd20529;
    data[16044] =  'sd20138;
    data[16045] = -'sd22875;
    data[16046] =  'sd3716;
    data[16047] =  'sd26012;
    data[16048] =  'sd18243;
    data[16049] = -'sd36140;
    data[16050] =  'sd74702;
    data[16051] =  'sd31391;
    data[16052] =  'sd55896;
    data[16053] =  'sd63590;
    data[16054] = -'sd46393;
    data[16055] =  'sd2931;
    data[16056] =  'sd20517;
    data[16057] = -'sd20222;
    data[16058] =  'sd22287;
    data[16059] = -'sd7832;
    data[16060] = -'sd54824;
    data[16061] = -'sd56086;
    data[16062] = -'sd64920;
    data[16063] =  'sd37083;
    data[16064] = -'sd68101;
    data[16065] =  'sd14816;
    data[16066] = -'sd60129;
    data[16067] =  'sd70620;
    data[16068] =  'sd2817;
    data[16069] =  'sd19719;
    data[16070] = -'sd25808;
    data[16071] = -'sd16815;
    data[16072] =  'sd46136;
    data[16073] = -'sd4730;
    data[16074] = -'sd33110;
    data[16075] = -'sd67929;
    data[16076] =  'sd16020;
    data[16077] = -'sd51701;
    data[16078] = -'sd34225;
    data[16079] = -'sd75734;
    data[16080] = -'sd38615;
    data[16081] =  'sd57377;
    data[16082] =  'sd73957;
    data[16083] =  'sd26176;
    data[16084] =  'sd19391;
    data[16085] = -'sd28104;
    data[16086] = -'sd32887;
    data[16087] = -'sd66368;
    data[16088] =  'sd26947;
    data[16089] =  'sd24788;
    data[16090] =  'sd9675;
    data[16091] =  'sd67725;
    data[16092] = -'sd17448;
    data[16093] =  'sd41705;
    data[16094] = -'sd35747;
    data[16095] =  'sd77453;
    data[16096] =  'sd50648;
    data[16097] =  'sd26854;
    data[16098] =  'sd24137;
    data[16099] =  'sd5118;
    data[16100] =  'sd35826;
    data[16101] = -'sd76900;
    data[16102] = -'sd46777;
    data[16103] =  'sd243;
    data[16104] =  'sd1701;
    data[16105] =  'sd11907;
    data[16106] = -'sd80492;
    data[16107] = -'sd71921;
    data[16108] = -'sd11924;
    data[16109] =  'sd80373;
    data[16110] =  'sd71088;
    data[16111] =  'sd6093;
    data[16112] =  'sd42651;
    data[16113] = -'sd29125;
    data[16114] = -'sd40034;
    data[16115] =  'sd47444;
    data[16116] =  'sd4426;
    data[16117] =  'sd30982;
    data[16118] =  'sd53033;
    data[16119] =  'sd43549;
    data[16120] = -'sd22839;
    data[16121] =  'sd3968;
    data[16122] =  'sd27776;
    data[16123] =  'sd30591;
    data[16124] =  'sd50296;
    data[16125] =  'sd24390;
    data[16126] =  'sd6889;
    data[16127] =  'sd48223;
    data[16128] =  'sd9879;
    data[16129] =  'sd69153;
    data[16130] = -'sd7452;
    data[16131] = -'sd52164;
    data[16132] = -'sd37466;
    data[16133] =  'sd65420;
    data[16134] = -'sd33583;
    data[16135] = -'sd71240;
    data[16136] = -'sd7157;
    data[16137] = -'sd50099;
    data[16138] = -'sd23011;
    data[16139] =  'sd2764;
    data[16140] =  'sd19348;
    data[16141] = -'sd28405;
    data[16142] = -'sd34994;
    data[16143] = -'sd81117;
    data[16144] = -'sd76296;
    data[16145] = -'sd42549;
    data[16146] =  'sd29839;
    data[16147] =  'sd45032;
    data[16148] = -'sd12458;
    data[16149] =  'sd76635;
    data[16150] =  'sd44922;
    data[16151] = -'sd13228;
    data[16152] =  'sd71245;
    data[16153] =  'sd7192;
    data[16154] =  'sd50344;
    data[16155] =  'sd24726;
    data[16156] =  'sd9241;
    data[16157] =  'sd64687;
    data[16158] = -'sd38714;
    data[16159] =  'sd56684;
    data[16160] =  'sd69106;
    data[16161] = -'sd7781;
    data[16162] = -'sd54467;
    data[16163] = -'sd53587;
    data[16164] = -'sd47427;
    data[16165] = -'sd4307;
    data[16166] = -'sd30149;
    data[16167] = -'sd47202;
    data[16168] = -'sd2732;
    data[16169] = -'sd19124;
    data[16170] =  'sd29973;
    data[16171] =  'sd45970;
    data[16172] = -'sd5892;
    data[16173] = -'sd41244;
    data[16174] =  'sd38974;
    data[16175] = -'sd54864;
    data[16176] = -'sd56366;
    data[16177] = -'sd66880;
    data[16178] =  'sd23363;
    data[16179] = -'sd300;
    data[16180] = -'sd2100;
    data[16181] = -'sd14700;
    data[16182] =  'sd60941;
    data[16183] = -'sd64936;
    data[16184] =  'sd36971;
    data[16185] = -'sd68885;
    data[16186] =  'sd9328;
    data[16187] =  'sd65296;
    data[16188] = -'sd34451;
    data[16189] = -'sd77316;
    data[16190] = -'sd49689;
    data[16191] = -'sd20141;
    data[16192] =  'sd22854;
    data[16193] = -'sd3863;
    data[16194] = -'sd27041;
    data[16195] = -'sd25446;
    data[16196] = -'sd14281;
    data[16197] =  'sd63874;
    data[16198] = -'sd44405;
    data[16199] =  'sd16847;
    data[16200] = -'sd45912;
    data[16201] =  'sd6298;
    data[16202] =  'sd44086;
    data[16203] = -'sd19080;
    data[16204] =  'sd30281;
    data[16205] =  'sd48126;
    data[16206] =  'sd9200;
    data[16207] =  'sd64400;
    data[16208] = -'sd40723;
    data[16209] =  'sd42621;
    data[16210] = -'sd29335;
    data[16211] = -'sd41504;
    data[16212] =  'sd37154;
    data[16213] = -'sd67604;
    data[16214] =  'sd18295;
    data[16215] = -'sd35776;
    data[16216] =  'sd77250;
    data[16217] =  'sd49227;
    data[16218] =  'sd16907;
    data[16219] = -'sd45492;
    data[16220] =  'sd9238;
    data[16221] =  'sd64666;
    data[16222] = -'sd38861;
    data[16223] =  'sd55655;
    data[16224] =  'sd61903;
    data[16225] = -'sd58202;
    data[16226] = -'sd79732;
    data[16227] = -'sd66601;
    data[16228] =  'sd25316;
    data[16229] =  'sd13371;
    data[16230] = -'sd70244;
    data[16231] = -'sd185;
    data[16232] = -'sd1295;
    data[16233] = -'sd9065;
    data[16234] = -'sd63455;
    data[16235] =  'sd47338;
    data[16236] =  'sd3684;
    data[16237] =  'sd25788;
    data[16238] =  'sd16675;
    data[16239] = -'sd47116;
    data[16240] = -'sd2130;
    data[16241] = -'sd14910;
    data[16242] =  'sd59471;
    data[16243] = -'sd75226;
    data[16244] = -'sd35059;
    data[16245] = -'sd81572;
    data[16246] = -'sd79481;
    data[16247] = -'sd64844;
    data[16248] =  'sd37615;
    data[16249] = -'sd64377;
    data[16250] =  'sd40884;
    data[16251] = -'sd41494;
    data[16252] =  'sd37224;
    data[16253] = -'sd67114;
    data[16254] =  'sd21725;
    data[16255] = -'sd11766;
    data[16256] =  'sd81479;
    data[16257] =  'sd78830;
    data[16258] =  'sd60287;
    data[16259] = -'sd69514;
    data[16260] =  'sd4925;
    data[16261] =  'sd34475;
    data[16262] =  'sd77484;
    data[16263] =  'sd50865;
    data[16264] =  'sd28373;
    data[16265] =  'sd34770;
    data[16266] =  'sd79549;
    data[16267] =  'sd65320;
    data[16268] = -'sd34283;
    data[16269] = -'sd76140;
    data[16270] = -'sd41457;
    data[16271] =  'sd37483;
    data[16272] = -'sd65301;
    data[16273] =  'sd34416;
    data[16274] =  'sd77071;
    data[16275] =  'sd47974;
    data[16276] =  'sd8136;
    data[16277] =  'sd56952;
    data[16278] =  'sd70982;
    data[16279] =  'sd5351;
    data[16280] =  'sd37457;
    data[16281] = -'sd65483;
    data[16282] =  'sd33142;
    data[16283] =  'sd68153;
    data[16284] = -'sd14452;
    data[16285] =  'sd62677;
    data[16286] = -'sd52784;
    data[16287] = -'sd41806;
    data[16288] =  'sd35040;
    data[16289] =  'sd81439;
    data[16290] =  'sd78550;
    data[16291] =  'sd58327;
    data[16292] =  'sd80607;
    data[16293] =  'sd72726;
    data[16294] =  'sd17559;
    data[16295] = -'sd40928;
    data[16296] =  'sd41186;
    data[16297] = -'sd39380;
    data[16298] =  'sd52022;
    data[16299] =  'sd36472;
    data[16300] = -'sd72378;
    data[16301] = -'sd15123;
    data[16302] =  'sd57980;
    data[16303] =  'sd78178;
    data[16304] =  'sd55723;
    data[16305] =  'sd62379;
    data[16306] = -'sd54870;
    data[16307] = -'sd56408;
    data[16308] = -'sd67174;
    data[16309] =  'sd21305;
    data[16310] = -'sd14706;
    data[16311] =  'sd60899;
    data[16312] = -'sd65230;
    data[16313] =  'sd34913;
    data[16314] =  'sd80550;
    data[16315] =  'sd72327;
    data[16316] =  'sd14766;
    data[16317] = -'sd60479;
    data[16318] =  'sd68170;
    data[16319] = -'sd14333;
    data[16320] =  'sd63510;
    data[16321] = -'sd46953;
    data[16322] = -'sd989;
    data[16323] = -'sd6923;
    data[16324] = -'sd48461;
    data[16325] = -'sd11545;
    data[16326] = -'sd80815;
    data[16327] = -'sd74182;
    data[16328] = -'sd27751;
    data[16329] = -'sd30416;
    data[16330] = -'sd49071;
    data[16331] = -'sd15815;
    data[16332] =  'sd53136;
    data[16333] =  'sd44270;
    data[16334] = -'sd17792;
    data[16335] =  'sd39297;
    data[16336] = -'sd52603;
    data[16337] = -'sd40539;
    data[16338] =  'sd43909;
    data[16339] = -'sd20319;
    data[16340] =  'sd21608;
    data[16341] = -'sd12585;
    data[16342] =  'sd75746;
    data[16343] =  'sd38699;
    data[16344] = -'sd56789;
    data[16345] = -'sd69841;
    data[16346] =  'sd2636;
    data[16347] =  'sd18452;
    data[16348] = -'sd34677;
    data[16349] = -'sd78898;
    data[16350] = -'sd60763;
    data[16351] =  'sd66182;
    data[16352] = -'sd28249;
    data[16353] = -'sd33902;
    data[16354] = -'sd73473;
    data[16355] = -'sd22788;
    data[16356] =  'sd4325;
    data[16357] =  'sd30275;
    data[16358] =  'sd48084;
    data[16359] =  'sd8906;
    data[16360] =  'sd62342;
    data[16361] = -'sd55129;
    data[16362] = -'sd58221;
    data[16363] = -'sd79865;
    data[16364] = -'sd67532;
    data[16365] =  'sd18799;
    data[16366] = -'sd32248;
    data[16367] = -'sd61895;
    data[16368] =  'sd58258;
    data[16369] =  'sd80124;
    data[16370] =  'sd69345;
    data[16371] = -'sd6108;
    data[16372] = -'sd42756;
    data[16373] =  'sd28390;
    data[16374] =  'sd34889;
    data[16375] =  'sd80382;
    data[16376] =  'sd71151;
    data[16377] =  'sd6534;
    data[16378] =  'sd45738;
    data[16379] = -'sd7516;
    data[16380] = -'sd52612;
    data[16381] = -'sd40602;
    data[16382] =  'sd43468;
    data[16383] = -'sd23406;
  end

endmodule

