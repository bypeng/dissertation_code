module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd761;
  localparam R_DEPTH = 'd10;
  localparam B_LEN = 'd1007;
  localparam B_DEPTH = 'd10;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [13: 0] in_data;
  input      [ 9: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 14'h004d; // 'd77
      10'd1    : in_data <= 14'h00f5; // 'd245
      10'd2    : in_data <= 14'h0068; // 'd104
      10'd3    : in_data <= 14'h02b1; // 'd689
      10'd4    : in_data <= 14'h0345; // 'd837
      10'd5    : in_data <= 14'h0406; // 'd1030
      10'd6    : in_data <= 14'h00e6; // 'd230
      10'd7    : in_data <= 14'h0337; // 'd823
      10'd8    : in_data <= 14'h05c3; // 'd1475
      10'd9    : in_data <= 14'h0472; // 'd1138
      10'd10   : in_data <= 14'h0202; // 'd514
      10'd11   : in_data <= 14'h00c5; // 'd197
      10'd12   : in_data <= 14'h04d2; // 'd1234
      10'd13   : in_data <= 14'h04c3; // 'd1219
      10'd14   : in_data <= 14'h0058; // 'd88
      10'd15   : in_data <= 14'h00f2; // 'd242
      10'd16   : in_data <= 14'h034e; // 'd846
      10'd17   : in_data <= 14'h05de; // 'd1502
      10'd18   : in_data <= 14'h0031; // 'd49
      10'd19   : in_data <= 14'h0196; // 'd406
      10'd20   : in_data <= 14'h04fc; // 'd1276
      10'd21   : in_data <= 14'h021e; // 'd542
      10'd22   : in_data <= 14'h0033; // 'd51
      10'd23   : in_data <= 14'h02e8; // 'd744
      10'd24   : in_data <= 14'h0080; // 'd128
      10'd25   : in_data <= 14'h029b; // 'd667
      10'd26   : in_data <= 14'h0054; // 'd84
      10'd27   : in_data <= 14'h0162; // 'd354
      10'd28   : in_data <= 14'h0046; // 'd70
      10'd29   : in_data <= 14'h01f0; // 'd496
      10'd30   : in_data <= 14'h040f; // 'd1039
      10'd31   : in_data <= 14'h05d5; // 'd1493
      10'd32   : in_data <= 14'h0380; // 'd896
      10'd33   : in_data <= 14'h0524; // 'd1316
      10'd34   : in_data <= 14'h00ec; // 'd236
      10'd35   : in_data <= 14'h038e; // 'd910
      10'd36   : in_data <= 14'h0072; // 'd114
      10'd37   : in_data <= 14'h0496; // 'd1174
      10'd38   : in_data <= 14'h0150; // 'd336
      10'd39   : in_data <= 14'h01cc; // 'd460
      10'd40   : in_data <= 14'h024a; // 'd586
      10'd41   : in_data <= 14'h05b1; // 'd1457
      10'd42   : in_data <= 14'h0360; // 'd864
      10'd43   : in_data <= 14'h0057; // 'd87
      10'd44   : in_data <= 14'h03f0; // 'd1008
      10'd45   : in_data <= 14'h0347; // 'd839
      10'd46   : in_data <= 14'h037f; // 'd895
      10'd47   : in_data <= 14'h05b2; // 'd1458
      10'd48   : in_data <= 14'h00ff; // 'd255
      10'd49   : in_data <= 14'h0526; // 'd1318
      10'd50   : in_data <= 14'h0018; // 'd24
      10'd51   : in_data <= 14'h01cf; // 'd463
      10'd52   : in_data <= 14'h0314; // 'd788
      10'd53   : in_data <= 14'h005e; // 'd94
      10'd54   : in_data <= 14'h02ff; // 'd767
      10'd55   : in_data <= 14'h0215; // 'd533
      10'd56   : in_data <= 14'h02b0; // 'd688
      10'd57   : in_data <= 14'h03d1; // 'd977
      10'd58   : in_data <= 14'h0250; // 'd592
      10'd59   : in_data <= 14'h02c7; // 'd711
      10'd60   : in_data <= 14'h01e0; // 'd480
      10'd61   : in_data <= 14'h0526; // 'd1318
      10'd62   : in_data <= 14'h02bb; // 'd699
      10'd63   : in_data <= 14'h0170; // 'd368
      10'd64   : in_data <= 14'h0423; // 'd1059
      10'd65   : in_data <= 14'h018b; // 'd395
      10'd66   : in_data <= 14'h0283; // 'd643
      10'd67   : in_data <= 14'h031e; // 'd798
      10'd68   : in_data <= 14'h0076; // 'd118
      10'd69   : in_data <= 14'h0042; // 'd66
      10'd70   : in_data <= 14'h01de; // 'd478
      10'd71   : in_data <= 14'h04d4; // 'd1236
      10'd72   : in_data <= 14'h04ba; // 'd1210
      10'd73   : in_data <= 14'h02c7; // 'd711
      10'd74   : in_data <= 14'h05c1; // 'd1473
      10'd75   : in_data <= 14'h059b; // 'd1435
      10'd76   : in_data <= 14'h0498; // 'd1176
      10'd77   : in_data <= 14'h0161; // 'd353
      10'd78   : in_data <= 14'h0379; // 'd889
      10'd79   : in_data <= 14'h03c1; // 'd961
      10'd80   : in_data <= 14'h002d; // 'd45
      10'd81   : in_data <= 14'h017e; // 'd382
      10'd82   : in_data <= 14'h043f; // 'd1087
      10'd83   : in_data <= 14'h03dd; // 'd989
      10'd84   : in_data <= 14'h01b3; // 'd435
      10'd85   : in_data <= 14'h0016; // 'd22
      10'd86   : in_data <= 14'h01ab; // 'd427
      10'd87   : in_data <= 14'h04e4; // 'd1252
      10'd88   : in_data <= 14'h04c4; // 'd1220
      10'd89   : in_data <= 14'h0519; // 'd1305
      10'd90   : in_data <= 14'h0585; // 'd1413
      10'd91   : in_data <= 14'h058a; // 'd1418
      10'd92   : in_data <= 14'h0115; // 'd277
      10'd93   : in_data <= 14'h02fa; // 'd762
      10'd94   : in_data <= 14'h03e7; // 'd999
      10'd95   : in_data <= 14'h02c2; // 'd706
      10'd96   : in_data <= 14'h014b; // 'd331
      10'd97   : in_data <= 14'h0568; // 'd1384
      10'd98   : in_data <= 14'h05f4; // 'd1524
      10'd99   : in_data <= 14'h04da; // 'd1242
      10'd100  : in_data <= 14'h01ab; // 'd427
      10'd101  : in_data <= 14'h0183; // 'd387
      10'd102  : in_data <= 14'h04c1; // 'd1217
      10'd103  : in_data <= 14'h0463; // 'd1123
      10'd104  : in_data <= 14'h01d2; // 'd466
      10'd105  : in_data <= 14'h002e; // 'd46
      10'd106  : in_data <= 14'h04f2; // 'd1266
      10'd107  : in_data <= 14'h00a3; // 'd163
      10'd108  : in_data <= 14'h05c0; // 'd1472
      10'd109  : in_data <= 14'h00cd; // 'd205
      10'd110  : in_data <= 14'h03bb; // 'd955
      10'd111  : in_data <= 14'h00ae; // 'd174
      10'd112  : in_data <= 14'h0023; // 'd35
      10'd113  : in_data <= 14'h02ee; // 'd750
      10'd114  : in_data <= 14'h055e; // 'd1374
      10'd115  : in_data <= 14'h0531; // 'd1329
      10'd116  : in_data <= 14'h047e; // 'd1150
      10'd117  : in_data <= 14'h02d0; // 'd720
      10'd118  : in_data <= 14'h0559; // 'd1369
      10'd119  : in_data <= 14'h02f8; // 'd760
      10'd120  : in_data <= 14'h02ad; // 'd685
      10'd121  : in_data <= 14'h053e; // 'd1342
      10'd122  : in_data <= 14'h001a; // 'd26
      10'd123  : in_data <= 14'h002c; // 'd44
      10'd124  : in_data <= 14'h00ba; // 'd186
      10'd125  : in_data <= 14'h05c4; // 'd1476
      10'd126  : in_data <= 14'h04d1; // 'd1233
      10'd127  : in_data <= 14'h010a; // 'd266
      10'd128  : in_data <= 14'h0173; // 'd371
      10'd129  : in_data <= 14'h01cf; // 'd463
      10'd130  : in_data <= 14'h056f; // 'd1391
      10'd131  : in_data <= 14'h0130; // 'd304
      10'd132  : in_data <= 14'h0103; // 'd259
      10'd133  : in_data <= 14'h043a; // 'd1082
      10'd134  : in_data <= 14'h00f3; // 'd243
      10'd135  : in_data <= 14'h0299; // 'd665
      10'd136  : in_data <= 14'h0095; // 'd149
      10'd137  : in_data <= 14'h034b; // 'd843
      10'd138  : in_data <= 14'h041e; // 'd1054
      10'd139  : in_data <= 14'h01bf; // 'd447
      10'd140  : in_data <= 14'h02dc; // 'd732
      10'd141  : in_data <= 14'h0348; // 'd840
      10'd142  : in_data <= 14'h0082; // 'd130
      10'd143  : in_data <= 14'h0478; // 'd1144
      10'd144  : in_data <= 14'h035b; // 'd859
      10'd145  : in_data <= 14'h017a; // 'd378
      10'd146  : in_data <= 14'h0231; // 'd561
      10'd147  : in_data <= 14'h0006; // 'd6
      10'd148  : in_data <= 14'h05d8; // 'd1496
      10'd149  : in_data <= 14'h0471; // 'd1137
      10'd150  : in_data <= 14'h0311; // 'd785
      10'd151  : in_data <= 14'h0159; // 'd345
      10'd152  : in_data <= 14'h0091; // 'd145
      10'd153  : in_data <= 14'h00e5; // 'd229
      10'd154  : in_data <= 14'h052b; // 'd1323
      10'd155  : in_data <= 14'h02c4; // 'd708
      10'd156  : in_data <= 14'h03b3; // 'd947
      10'd157  : in_data <= 14'h0113; // 'd275
      10'd158  : in_data <= 14'h014d; // 'd333
      10'd159  : in_data <= 14'h002e; // 'd46
      10'd160  : in_data <= 14'h0445; // 'd1093
      10'd161  : in_data <= 14'h02a4; // 'd676
      10'd162  : in_data <= 14'h0217; // 'd535
      10'd163  : in_data <= 14'h00b7; // 'd183
      10'd164  : in_data <= 14'h00de; // 'd222
      10'd165  : in_data <= 14'h0491; // 'd1169
      10'd166  : in_data <= 14'h00d3; // 'd211
      10'd167  : in_data <= 14'h0033; // 'd51
      10'd168  : in_data <= 14'h0237; // 'd567
      10'd169  : in_data <= 14'h03d8; // 'd984
      10'd170  : in_data <= 14'h03bc; // 'd956
      10'd171  : in_data <= 14'h022d; // 'd557
      10'd172  : in_data <= 14'h0511; // 'd1297
      10'd173  : in_data <= 14'h05ab; // 'd1451
      10'd174  : in_data <= 14'h0521; // 'd1313
      10'd175  : in_data <= 14'h02ac; // 'd684
      10'd176  : in_data <= 14'h05f7; // 'd1527
      10'd177  : in_data <= 14'h0109; // 'd265
      10'd178  : in_data <= 14'h013e; // 'd318
      10'd179  : in_data <= 14'h03d8; // 'd984
      10'd180  : in_data <= 14'h006e; // 'd110
      10'd181  : in_data <= 14'h050d; // 'd1293
      10'd182  : in_data <= 14'h0132; // 'd306
      10'd183  : in_data <= 14'h00d7; // 'd215
      10'd184  : in_data <= 14'h0309; // 'd777
      10'd185  : in_data <= 14'h02c2; // 'd706
      10'd186  : in_data <= 14'h03bb; // 'd955
      10'd187  : in_data <= 14'h048b; // 'd1163
      10'd188  : in_data <= 14'h02b6; // 'd694
      10'd189  : in_data <= 14'h0293; // 'd659
      10'd190  : in_data <= 14'h045e; // 'd1118
      10'd191  : in_data <= 14'h0099; // 'd153
      10'd192  : in_data <= 14'h0014; // 'd20
      10'd193  : in_data <= 14'h00c0; // 'd192
      10'd194  : in_data <= 14'h02ba; // 'd698
      10'd195  : in_data <= 14'h0595; // 'd1429
      10'd196  : in_data <= 14'h01f8; // 'd504
      10'd197  : in_data <= 14'h05b2; // 'd1458
      10'd198  : in_data <= 14'h0334; // 'd820
      10'd199  : in_data <= 14'h037d; // 'd893
      10'd200  : in_data <= 14'h0102; // 'd258
      10'd201  : in_data <= 14'h01c0; // 'd448
      10'd202  : in_data <= 14'h03cf; // 'd975
      10'd203  : in_data <= 14'h0359; // 'd857
      10'd204  : in_data <= 14'h00ae; // 'd174
      10'd205  : in_data <= 14'h0090; // 'd144
      10'd206  : in_data <= 14'h01e4; // 'd484
      10'd207  : in_data <= 14'h00a1; // 'd161
      10'd208  : in_data <= 14'h011e; // 'd286
      10'd209  : in_data <= 14'h0144; // 'd324
      10'd210  : in_data <= 14'h0212; // 'd530
      10'd211  : in_data <= 14'h014c; // 'd332
      10'd212  : in_data <= 14'h03a6; // 'd934
      10'd213  : in_data <= 14'h003c; // 'd60
      10'd214  : in_data <= 14'h037f; // 'd895
      10'd215  : in_data <= 14'h0396; // 'd918
      10'd216  : in_data <= 14'h039f; // 'd927
      10'd217  : in_data <= 14'h02bf; // 'd703
      10'd218  : in_data <= 14'h05f0; // 'd1520
      10'd219  : in_data <= 14'h0583; // 'd1411
      10'd220  : in_data <= 14'h0319; // 'd793
      10'd221  : in_data <= 14'h053a; // 'd1338
      10'd222  : in_data <= 14'h0251; // 'd593
      10'd223  : in_data <= 14'h02d2; // 'd722
      10'd224  : in_data <= 14'h05be; // 'd1470
      10'd225  : in_data <= 14'h00d8; // 'd216
      10'd226  : in_data <= 14'h0594; // 'd1428
      10'd227  : in_data <= 14'h02bf; // 'd703
      10'd228  : in_data <= 14'h008c; // 'd140
      10'd229  : in_data <= 14'h03a7; // 'd935
      10'd230  : in_data <= 14'h0083; // 'd131
      10'd231  : in_data <= 14'h0089; // 'd137
      10'd232  : in_data <= 14'h0214; // 'd532
      10'd233  : in_data <= 14'h01af; // 'd431
      10'd234  : in_data <= 14'h05c0; // 'd1472
      10'd235  : in_data <= 14'h0242; // 'd578
      10'd236  : in_data <= 14'h01fd; // 'd509
      10'd237  : in_data <= 14'h02bc; // 'd700
      10'd238  : in_data <= 14'h0107; // 'd263
      10'd239  : in_data <= 14'h045b; // 'd1115
      10'd240  : in_data <= 14'h0179; // 'd377
      10'd241  : in_data <= 14'h02c0; // 'd704
      10'd242  : in_data <= 14'h05f4; // 'd1524
      10'd243  : in_data <= 14'h0438; // 'd1080
      10'd244  : in_data <= 14'h014e; // 'd334
      10'd245  : in_data <= 14'h035e; // 'd862
      10'd246  : in_data <= 14'h0038; // 'd56
      10'd247  : in_data <= 14'h0563; // 'd1379
      10'd248  : in_data <= 14'h0024; // 'd36
      10'd249  : in_data <= 14'h008d; // 'd141
      10'd250  : in_data <= 14'h00a2; // 'd162
      10'd251  : in_data <= 14'h0568; // 'd1384
      10'd252  : in_data <= 14'h037f; // 'd895
      10'd253  : in_data <= 14'h010b; // 'd267
      10'd254  : in_data <= 14'h053e; // 'd1342
      10'd255  : in_data <= 14'h02f6; // 'd758
      10'd256  : in_data <= 14'h05c7; // 'd1479
      10'd257  : in_data <= 14'h02e3; // 'd739
      10'd258  : in_data <= 14'h0074; // 'd116
      10'd259  : in_data <= 14'h0180; // 'd384
      10'd260  : in_data <= 14'h0044; // 'd68
      10'd261  : in_data <= 14'h01fb; // 'd507
      10'd262  : in_data <= 14'h01bc; // 'd444
      10'd263  : in_data <= 14'h01fa; // 'd506
      10'd264  : in_data <= 14'h0270; // 'd624
      10'd265  : in_data <= 14'h0593; // 'd1427
      10'd266  : in_data <= 14'h025b; // 'd603
      10'd267  : in_data <= 14'h018e; // 'd398
      10'd268  : in_data <= 14'h05a6; // 'd1446
      10'd269  : in_data <= 14'h0370; // 'd880
      10'd270  : in_data <= 14'h03dc; // 'd988
      10'd271  : in_data <= 14'h02f7; // 'd759
      10'd272  : in_data <= 14'h00ce; // 'd206
      10'd273  : in_data <= 14'h038d; // 'd909
      10'd274  : in_data <= 14'h02ea; // 'd746
      10'd275  : in_data <= 14'h00f1; // 'd241
      10'd276  : in_data <= 14'h00a3; // 'd163
      10'd277  : in_data <= 14'h008c; // 'd140
      10'd278  : in_data <= 14'h0282; // 'd642
      10'd279  : in_data <= 14'h0233; // 'd563
      10'd280  : in_data <= 14'h03b3; // 'd947
      10'd281  : in_data <= 14'h04d7; // 'd1239
      10'd282  : in_data <= 14'h025d; // 'd605
      10'd283  : in_data <= 14'h046a; // 'd1130
      10'd284  : in_data <= 14'h0410; // 'd1040
      10'd285  : in_data <= 14'h0115; // 'd277
      10'd286  : in_data <= 14'h01ac; // 'd428
      10'd287  : in_data <= 14'h0564; // 'd1380
      10'd288  : in_data <= 14'h00f5; // 'd245
      10'd289  : in_data <= 14'h04da; // 'd1242
      10'd290  : in_data <= 14'h00d6; // 'd214
      10'd291  : in_data <= 14'h051f; // 'd1311
      10'd292  : in_data <= 14'h023f; // 'd575
      10'd293  : in_data <= 14'h04c7; // 'd1223
      10'd294  : in_data <= 14'h040a; // 'd1034
      10'd295  : in_data <= 14'h0320; // 'd800
      10'd296  : in_data <= 14'h04e8; // 'd1256
      10'd297  : in_data <= 14'h04ac; // 'd1196
      10'd298  : in_data <= 14'h04dd; // 'd1245
      10'd299  : in_data <= 14'h04f3; // 'd1267
      10'd300  : in_data <= 14'h01d6; // 'd470
      10'd301  : in_data <= 14'h039f; // 'd927
      10'd302  : in_data <= 14'h0405; // 'd1029
      10'd303  : in_data <= 14'h01b5; // 'd437
      10'd304  : in_data <= 14'h03d9; // 'd985
      10'd305  : in_data <= 14'h0520; // 'd1312
      10'd306  : in_data <= 14'h014f; // 'd335
      10'd307  : in_data <= 14'h0313; // 'd787
      10'd308  : in_data <= 14'h0073; // 'd115
      10'd309  : in_data <= 14'h033d; // 'd829
      10'd310  : in_data <= 14'h04ea; // 'd1258
      10'd311  : in_data <= 14'h034d; // 'd845
      10'd312  : in_data <= 14'h013e; // 'd318
      10'd313  : in_data <= 14'h042a; // 'd1066
      10'd314  : in_data <= 14'h0346; // 'd838
      10'd315  : in_data <= 14'h03a9; // 'd937
      10'd316  : in_data <= 14'h01a5; // 'd421
      10'd317  : in_data <= 14'h0057; // 'd87
      10'd318  : in_data <= 14'h041a; // 'd1050
      10'd319  : in_data <= 14'h0414; // 'd1044
      10'd320  : in_data <= 14'h00aa; // 'd170
      10'd321  : in_data <= 14'h054e; // 'd1358
      10'd322  : in_data <= 14'h005d; // 'd93
      10'd323  : in_data <= 14'h044f; // 'd1103
      10'd324  : in_data <= 14'h021e; // 'd542
      10'd325  : in_data <= 14'h04f0; // 'd1264
      10'd326  : in_data <= 14'h00fa; // 'd250
      10'd327  : in_data <= 14'h0311; // 'd785
      10'd328  : in_data <= 14'h00b8; // 'd184
      10'd329  : in_data <= 14'h04fa; // 'd1274
      10'd330  : in_data <= 14'h03fa; // 'd1018
      10'd331  : in_data <= 14'h04d5; // 'd1237
      10'd332  : in_data <= 14'h05ae; // 'd1454
      10'd333  : in_data <= 14'h0389; // 'd905
      10'd334  : in_data <= 14'h01d3; // 'd467
      10'd335  : in_data <= 14'h054f; // 'd1359
      10'd336  : in_data <= 14'h0430; // 'd1072
      10'd337  : in_data <= 14'h03ea; // 'd1002
      10'd338  : in_data <= 14'h05e0; // 'd1504
      10'd339  : in_data <= 14'h038c; // 'd908
      10'd340  : in_data <= 14'h0010; // 'd16
      10'd341  : in_data <= 14'h0594; // 'd1428
      10'd342  : in_data <= 14'h03ba; // 'd954
      10'd343  : in_data <= 14'h05cb; // 'd1483
      10'd344  : in_data <= 14'h0459; // 'd1113
      10'd345  : in_data <= 14'h0468; // 'd1128
      10'd346  : in_data <= 14'h0309; // 'd777
      10'd347  : in_data <= 14'h01c7; // 'd455
      10'd348  : in_data <= 14'h004d; // 'd77
      10'd349  : in_data <= 14'h02b8; // 'd696
      10'd350  : in_data <= 14'h01da; // 'd474
      10'd351  : in_data <= 14'h047b; // 'd1147
      10'd352  : in_data <= 14'h00c9; // 'd201
      10'd353  : in_data <= 14'h010b; // 'd267
      10'd354  : in_data <= 14'h05d6; // 'd1494
      10'd355  : in_data <= 14'h040f; // 'd1039
      10'd356  : in_data <= 14'h006b; // 'd107
      10'd357  : in_data <= 14'h0300; // 'd768
      10'd358  : in_data <= 14'h0304; // 'd772
      10'd359  : in_data <= 14'h05e5; // 'd1509
      10'd360  : in_data <= 14'h04c1; // 'd1217
      10'd361  : in_data <= 14'h0028; // 'd40
      10'd362  : in_data <= 14'h057d; // 'd1405
      10'd363  : in_data <= 14'h0495; // 'd1173
      10'd364  : in_data <= 14'h00a1; // 'd161
      10'd365  : in_data <= 14'h0143; // 'd323
      10'd366  : in_data <= 14'h00a0; // 'd160
      10'd367  : in_data <= 14'h050b; // 'd1291
      10'd368  : in_data <= 14'h01dc; // 'd476
      10'd369  : in_data <= 14'h03a3; // 'd931
      10'd370  : in_data <= 14'h031c; // 'd796
      10'd371  : in_data <= 14'h0032; // 'd50
      10'd372  : in_data <= 14'h002c; // 'd44
      10'd373  : in_data <= 14'h0541; // 'd1345
      10'd374  : in_data <= 14'h00d2; // 'd210
      10'd375  : in_data <= 14'h0498; // 'd1176
      10'd376  : in_data <= 14'h0587; // 'd1415
      10'd377  : in_data <= 14'h056b; // 'd1387
      10'd378  : in_data <= 14'h05c1; // 'd1473
      10'd379  : in_data <= 14'h0031; // 'd49
      10'd380  : in_data <= 14'h03d3; // 'd979
      10'd381  : in_data <= 14'h046c; // 'd1132
      10'd382  : in_data <= 14'h00ea; // 'd234
      10'd383  : in_data <= 14'h0036; // 'd54
      10'd384  : in_data <= 14'h03f3; // 'd1011
      10'd385  : in_data <= 14'h008c; // 'd140
      10'd386  : in_data <= 14'h014c; // 'd332
      10'd387  : in_data <= 14'h0499; // 'd1177
      10'd388  : in_data <= 14'h05b2; // 'd1458
      10'd389  : in_data <= 14'h04d9; // 'd1241
      10'd390  : in_data <= 14'h051c; // 'd1308
      10'd391  : in_data <= 14'h0258; // 'd600
      10'd392  : in_data <= 14'h04fd; // 'd1277
      10'd393  : in_data <= 14'h0394; // 'd916
      10'd394  : in_data <= 14'h0181; // 'd385
      10'd395  : in_data <= 14'h0435; // 'd1077
      10'd396  : in_data <= 14'h029b; // 'd667
      10'd397  : in_data <= 14'h038e; // 'd910
      10'd398  : in_data <= 14'h03cf; // 'd975
      10'd399  : in_data <= 14'h05c5; // 'd1477
      10'd400  : in_data <= 14'h057f; // 'd1407
      10'd401  : in_data <= 14'h0522; // 'd1314
      10'd402  : in_data <= 14'h05cf; // 'd1487
      10'd403  : in_data <= 14'h0392; // 'd914
      10'd404  : in_data <= 14'h00ac; // 'd172
      10'd405  : in_data <= 14'h007c; // 'd124
      10'd406  : in_data <= 14'h00bb; // 'd187
      10'd407  : in_data <= 14'h05d2; // 'd1490
      10'd408  : in_data <= 14'h03b8; // 'd952
      10'd409  : in_data <= 14'h03ba; // 'd954
      10'd410  : in_data <= 14'h03d2; // 'd978
      10'd411  : in_data <= 14'h00a4; // 'd164
      10'd412  : in_data <= 14'h03e9; // 'd1001
      10'd413  : in_data <= 14'h03a5; // 'd933
      10'd414  : in_data <= 14'h0167; // 'd359
      10'd415  : in_data <= 14'h01c3; // 'd451
      10'd416  : in_data <= 14'h02b1; // 'd689
      10'd417  : in_data <= 14'h0312; // 'd786
      10'd418  : in_data <= 14'h03cc; // 'd972
      10'd419  : in_data <= 14'h055a; // 'd1370
      10'd420  : in_data <= 14'h000b; // 'd11
      10'd421  : in_data <= 14'h0583; // 'd1411
      10'd422  : in_data <= 14'h0334; // 'd820
      10'd423  : in_data <= 14'h020b; // 'd523
      10'd424  : in_data <= 14'h0307; // 'd775
      10'd425  : in_data <= 14'h02ba; // 'd698
      10'd426  : in_data <= 14'h01c6; // 'd454
      10'd427  : in_data <= 14'h0199; // 'd409
      10'd428  : in_data <= 14'h0071; // 'd113
      10'd429  : in_data <= 14'h01dc; // 'd476
      10'd430  : in_data <= 14'h007f; // 'd127
      10'd431  : in_data <= 14'h0167; // 'd359
      10'd432  : in_data <= 14'h0429; // 'd1065
      10'd433  : in_data <= 14'h03f9; // 'd1017
      10'd434  : in_data <= 14'h02ce; // 'd718
      10'd435  : in_data <= 14'h02f1; // 'd753
      10'd436  : in_data <= 14'h01c0; // 'd448
      10'd437  : in_data <= 14'h03dd; // 'd989
      10'd438  : in_data <= 14'h01b7; // 'd439
      10'd439  : in_data <= 14'h02b1; // 'd689
      10'd440  : in_data <= 14'h00dc; // 'd220
      10'd441  : in_data <= 14'h009e; // 'd158
      10'd442  : in_data <= 14'h0224; // 'd548
      10'd443  : in_data <= 14'h0442; // 'd1090
      10'd444  : in_data <= 14'h04f1; // 'd1265
      10'd445  : in_data <= 14'h02ba; // 'd698
      10'd446  : in_data <= 14'h0033; // 'd51
      10'd447  : in_data <= 14'h0563; // 'd1379
      10'd448  : in_data <= 14'h025d; // 'd605
      10'd449  : in_data <= 14'h02cb; // 'd715
      10'd450  : in_data <= 14'h037b; // 'd891
      10'd451  : in_data <= 14'h0287; // 'd647
      10'd452  : in_data <= 14'h05de; // 'd1502
      10'd453  : in_data <= 14'h05c9; // 'd1481
      10'd454  : in_data <= 14'h0227; // 'd551
      10'd455  : in_data <= 14'h0569; // 'd1385
      10'd456  : in_data <= 14'h0463; // 'd1123
      10'd457  : in_data <= 14'h04dc; // 'd1244
      10'd458  : in_data <= 14'h04ba; // 'd1210
      10'd459  : in_data <= 14'h0164; // 'd356
      10'd460  : in_data <= 14'h027d; // 'd637
      10'd461  : in_data <= 14'h045e; // 'd1118
      10'd462  : in_data <= 14'h0530; // 'd1328
      10'd463  : in_data <= 14'h005e; // 'd94
      10'd464  : in_data <= 14'h057c; // 'd1404
      10'd465  : in_data <= 14'h052d; // 'd1325
      10'd466  : in_data <= 14'h033e; // 'd830
      10'd467  : in_data <= 14'h03ad; // 'd941
      10'd468  : in_data <= 14'h006f; // 'd111
      10'd469  : in_data <= 14'h00a2; // 'd162
      10'd470  : in_data <= 14'h00a9; // 'd169
      10'd471  : in_data <= 14'h0164; // 'd356
      10'd472  : in_data <= 14'h050c; // 'd1292
      10'd473  : in_data <= 14'h04e0; // 'd1248
      10'd474  : in_data <= 14'h01d1; // 'd465
      10'd475  : in_data <= 14'h0212; // 'd530
      10'd476  : in_data <= 14'h044f; // 'd1103
      10'd477  : in_data <= 14'h03bb; // 'd955
      10'd478  : in_data <= 14'h04e6; // 'd1254
      10'd479  : in_data <= 14'h04f0; // 'd1264
      10'd480  : in_data <= 14'h0318; // 'd792
      10'd481  : in_data <= 14'h04b9; // 'd1209
      10'd482  : in_data <= 14'h01e3; // 'd483
      10'd483  : in_data <= 14'h01c7; // 'd455
      10'd484  : in_data <= 14'h0542; // 'd1346
      10'd485  : in_data <= 14'h0194; // 'd404
      10'd486  : in_data <= 14'h0206; // 'd518
      10'd487  : in_data <= 14'h02a4; // 'd676
      10'd488  : in_data <= 14'h039a; // 'd922
      10'd489  : in_data <= 14'h03e5; // 'd997
      10'd490  : in_data <= 14'h04d5; // 'd1237
      10'd491  : in_data <= 14'h0084; // 'd132
      10'd492  : in_data <= 14'h009b; // 'd155
      10'd493  : in_data <= 14'h0297; // 'd663
      10'd494  : in_data <= 14'h01a0; // 'd416
      10'd495  : in_data <= 14'h0081; // 'd129
      10'd496  : in_data <= 14'h053e; // 'd1342
      10'd497  : in_data <= 14'h0221; // 'd545
      10'd498  : in_data <= 14'h02c7; // 'd711
      10'd499  : in_data <= 14'h0549; // 'd1353
      10'd500  : in_data <= 14'h052c; // 'd1324
      10'd501  : in_data <= 14'h0537; // 'd1335
      10'd502  : in_data <= 14'h0411; // 'd1041
      10'd503  : in_data <= 14'h0409; // 'd1033
      10'd504  : in_data <= 14'h0153; // 'd339
      10'd505  : in_data <= 14'h044b; // 'd1099
      10'd506  : in_data <= 14'h03e4; // 'd996
      10'd507  : in_data <= 14'h030e; // 'd782
      10'd508  : in_data <= 14'h006a; // 'd106
      10'd509  : in_data <= 14'h0267; // 'd615
      10'd510  : in_data <= 14'h0544; // 'd1348
      10'd511  : in_data <= 14'h03cd; // 'd973
      10'd512  : in_data <= 14'h01d6; // 'd470
      10'd513  : in_data <= 14'h013a; // 'd314
      10'd514  : in_data <= 14'h01d5; // 'd469
      10'd515  : in_data <= 14'h006d; // 'd109
      10'd516  : in_data <= 14'h01a0; // 'd416
      10'd517  : in_data <= 14'h00da; // 'd218
      10'd518  : in_data <= 14'h050f; // 'd1295
      10'd519  : in_data <= 14'h009c; // 'd156
      10'd520  : in_data <= 14'h00d0; // 'd208
      10'd521  : in_data <= 14'h05bb; // 'd1467
      10'd522  : in_data <= 14'h025b; // 'd603
      10'd523  : in_data <= 14'h01e4; // 'd484
      10'd524  : in_data <= 14'h0224; // 'd548
      10'd525  : in_data <= 14'h04b4; // 'd1204
      10'd526  : in_data <= 14'h04b2; // 'd1202
      10'd527  : in_data <= 14'h0321; // 'd801
      10'd528  : in_data <= 14'h0415; // 'd1045
      10'd529  : in_data <= 14'h005e; // 'd94
      10'd530  : in_data <= 14'h0589; // 'd1417
      10'd531  : in_data <= 14'h0250; // 'd592
      10'd532  : in_data <= 14'h05cd; // 'd1485
      10'd533  : in_data <= 14'h028d; // 'd653
      10'd534  : in_data <= 14'h03c5; // 'd965
      10'd535  : in_data <= 14'h010f; // 'd271
      10'd536  : in_data <= 14'h0509; // 'd1289
      10'd537  : in_data <= 14'h0218; // 'd536
      10'd538  : in_data <= 14'h025e; // 'd606
      10'd539  : in_data <= 14'h01fa; // 'd506
      10'd540  : in_data <= 14'h0139; // 'd313
      10'd541  : in_data <= 14'h0379; // 'd889
      10'd542  : in_data <= 14'h01a6; // 'd422
      10'd543  : in_data <= 14'h0002; // 'd2
      10'd544  : in_data <= 14'h0152; // 'd338
      10'd545  : in_data <= 14'h02ef; // 'd751
      10'd546  : in_data <= 14'h05c8; // 'd1480
      10'd547  : in_data <= 14'h0516; // 'd1302
      10'd548  : in_data <= 14'h04a2; // 'd1186
      10'd549  : in_data <= 14'h0016; // 'd22
      10'd550  : in_data <= 14'h0187; // 'd391
      10'd551  : in_data <= 14'h03e8; // 'd1000
      10'd552  : in_data <= 14'h040a; // 'd1034
      10'd553  : in_data <= 14'h0569; // 'd1385
      10'd554  : in_data <= 14'h0397; // 'd919
      10'd555  : in_data <= 14'h0126; // 'd294
      10'd556  : in_data <= 14'h04a5; // 'd1189
      10'd557  : in_data <= 14'h019a; // 'd410
      10'd558  : in_data <= 14'h0477; // 'd1143
      10'd559  : in_data <= 14'h05de; // 'd1502
      10'd560  : in_data <= 14'h021b; // 'd539
      10'd561  : in_data <= 14'h03ee; // 'd1006
      10'd562  : in_data <= 14'h0056; // 'd86
      10'd563  : in_data <= 14'h053f; // 'd1343
      10'd564  : in_data <= 14'h0224; // 'd548
      10'd565  : in_data <= 14'h0128; // 'd296
      10'd566  : in_data <= 14'h05d1; // 'd1489
      10'd567  : in_data <= 14'h050e; // 'd1294
      10'd568  : in_data <= 14'h048c; // 'd1164
      10'd569  : in_data <= 14'h057a; // 'd1402
      10'd570  : in_data <= 14'h0585; // 'd1413
      10'd571  : in_data <= 14'h035c; // 'd860
      10'd572  : in_data <= 14'h0244; // 'd580
      10'd573  : in_data <= 14'h0547; // 'd1351
      10'd574  : in_data <= 14'h043e; // 'd1086
      10'd575  : in_data <= 14'h0044; // 'd68
      10'd576  : in_data <= 14'h0109; // 'd265
      10'd577  : in_data <= 14'h04ce; // 'd1230
      10'd578  : in_data <= 14'h00be; // 'd190
      10'd579  : in_data <= 14'h04da; // 'd1242
      10'd580  : in_data <= 14'h00c5; // 'd197
      10'd581  : in_data <= 14'h005d; // 'd93
      10'd582  : in_data <= 14'h0437; // 'd1079
      10'd583  : in_data <= 14'h045f; // 'd1119
      10'd584  : in_data <= 14'h0502; // 'd1282
      10'd585  : in_data <= 14'h0566; // 'd1382
      10'd586  : in_data <= 14'h0377; // 'd887
      10'd587  : in_data <= 14'h0327; // 'd807
      10'd588  : in_data <= 14'h0350; // 'd848
      10'd589  : in_data <= 14'h01a6; // 'd422
      10'd590  : in_data <= 14'h01d9; // 'd473
      10'd591  : in_data <= 14'h0370; // 'd880
      10'd592  : in_data <= 14'h05f1; // 'd1521
      10'd593  : in_data <= 14'h034a; // 'd842
      10'd594  : in_data <= 14'h051c; // 'd1308
      10'd595  : in_data <= 14'h05c2; // 'd1474
      10'd596  : in_data <= 14'h05ba; // 'd1466
      10'd597  : in_data <= 14'h05f7; // 'd1527
      10'd598  : in_data <= 14'h03ee; // 'd1006
      10'd599  : in_data <= 14'h0008; // 'd8
      10'd600  : in_data <= 14'h0477; // 'd1143
      10'd601  : in_data <= 14'h03ed; // 'd1005
      10'd602  : in_data <= 14'h00f0; // 'd240
      10'd603  : in_data <= 14'h044f; // 'd1103
      10'd604  : in_data <= 14'h00bf; // 'd191
      10'd605  : in_data <= 14'h058b; // 'd1419
      10'd606  : in_data <= 14'h0186; // 'd390
      10'd607  : in_data <= 14'h040d; // 'd1037
      10'd608  : in_data <= 14'h02b2; // 'd690
      10'd609  : in_data <= 14'h0441; // 'd1089
      10'd610  : in_data <= 14'h042b; // 'd1067
      10'd611  : in_data <= 14'h0352; // 'd850
      10'd612  : in_data <= 14'h00ce; // 'd206
      10'd613  : in_data <= 14'h028b; // 'd651
      10'd614  : in_data <= 14'h021a; // 'd538
      10'd615  : in_data <= 14'h04b4; // 'd1204
      10'd616  : in_data <= 14'h00e3; // 'd227
      10'd617  : in_data <= 14'h005d; // 'd93
      10'd618  : in_data <= 14'h0003; // 'd3
      10'd619  : in_data <= 14'h03bc; // 'd956
      10'd620  : in_data <= 14'h0400; // 'd1024
      10'd621  : in_data <= 14'h02dc; // 'd732
      10'd622  : in_data <= 14'h0453; // 'd1107
      10'd623  : in_data <= 14'h0446; // 'd1094
      10'd624  : in_data <= 14'h025f; // 'd607
      10'd625  : in_data <= 14'h0244; // 'd580
      10'd626  : in_data <= 14'h00ec; // 'd236
      10'd627  : in_data <= 14'h05d7; // 'd1495
      10'd628  : in_data <= 14'h0059; // 'd89
      10'd629  : in_data <= 14'h0014; // 'd20
      10'd630  : in_data <= 14'h054c; // 'd1356
      10'd631  : in_data <= 14'h05dc; // 'd1500
      10'd632  : in_data <= 14'h03a3; // 'd931
      10'd633  : in_data <= 14'h02c1; // 'd705
      10'd634  : in_data <= 14'h055d; // 'd1373
      10'd635  : in_data <= 14'h00f4; // 'd244
      10'd636  : in_data <= 14'h05a4; // 'd1444
      10'd637  : in_data <= 14'h0196; // 'd406
      10'd638  : in_data <= 14'h01e5; // 'd485
      10'd639  : in_data <= 14'h0431; // 'd1073
      10'd640  : in_data <= 14'h0514; // 'd1300
      10'd641  : in_data <= 14'h0357; // 'd855
      10'd642  : in_data <= 14'h003b; // 'd59
      10'd643  : in_data <= 14'h0418; // 'd1048
      10'd644  : in_data <= 14'h013f; // 'd319
      10'd645  : in_data <= 14'h0128; // 'd296
      10'd646  : in_data <= 14'h043f; // 'd1087
      10'd647  : in_data <= 14'h03af; // 'd943
      10'd648  : in_data <= 14'h059a; // 'd1434
      10'd649  : in_data <= 14'h050f; // 'd1295
      10'd650  : in_data <= 14'h059e; // 'd1438
      10'd651  : in_data <= 14'h0411; // 'd1041
      10'd652  : in_data <= 14'h04a5; // 'd1189
      10'd653  : in_data <= 14'h03a8; // 'd936
      10'd654  : in_data <= 14'h0219; // 'd537
      10'd655  : in_data <= 14'h0288; // 'd648
      10'd656  : in_data <= 14'h02f7; // 'd759
      10'd657  : in_data <= 14'h00f9; // 'd249
      10'd658  : in_data <= 14'h024c; // 'd588
      10'd659  : in_data <= 14'h0152; // 'd338
      10'd660  : in_data <= 14'h01c2; // 'd450
      10'd661  : in_data <= 14'h0591; // 'd1425
      10'd662  : in_data <= 14'h0397; // 'd919
      10'd663  : in_data <= 14'h0145; // 'd325
      10'd664  : in_data <= 14'h0379; // 'd889
      10'd665  : in_data <= 14'h04fd; // 'd1277
      10'd666  : in_data <= 14'h0124; // 'd292
      10'd667  : in_data <= 14'h0078; // 'd120
      10'd668  : in_data <= 14'h019f; // 'd415
      10'd669  : in_data <= 14'h0056; // 'd86
      10'd670  : in_data <= 14'h01e9; // 'd489
      10'd671  : in_data <= 14'h01ec; // 'd492
      10'd672  : in_data <= 14'h0286; // 'd646
      10'd673  : in_data <= 14'h0051; // 'd81
      10'd674  : in_data <= 14'h0497; // 'd1175
      10'd675  : in_data <= 14'h05e8; // 'd1512
      10'd676  : in_data <= 14'h0317; // 'd791
      10'd677  : in_data <= 14'h004f; // 'd79
      10'd678  : in_data <= 14'h00ad; // 'd173
      10'd679  : in_data <= 14'h02a9; // 'd681
      10'd680  : in_data <= 14'h035f; // 'd863
      10'd681  : in_data <= 14'h02ba; // 'd698
      10'd682  : in_data <= 14'h0121; // 'd289
      10'd683  : in_data <= 14'h056d; // 'd1389
      10'd684  : in_data <= 14'h0222; // 'd546
      10'd685  : in_data <= 14'h0540; // 'd1344
      10'd686  : in_data <= 14'h0372; // 'd882
      10'd687  : in_data <= 14'h015e; // 'd350
      10'd688  : in_data <= 14'h001c; // 'd28
      10'd689  : in_data <= 14'h0074; // 'd116
      10'd690  : in_data <= 14'h0218; // 'd536
      10'd691  : in_data <= 14'h01c6; // 'd454
      10'd692  : in_data <= 14'h038e; // 'd910
      10'd693  : in_data <= 14'h0359; // 'd857
      10'd694  : in_data <= 14'h021a; // 'd538
      10'd695  : in_data <= 14'h01f2; // 'd498
      10'd696  : in_data <= 14'h059e; // 'd1438
      10'd697  : in_data <= 14'h0354; // 'd852
      10'd698  : in_data <= 14'h03e6; // 'd998
      10'd699  : in_data <= 14'h01cb; // 'd459
      10'd700  : in_data <= 14'h0495; // 'd1173
      10'd701  : in_data <= 14'h017c; // 'd380
      10'd702  : in_data <= 14'h0498; // 'd1176
      10'd703  : in_data <= 14'h0404; // 'd1028
      10'd704  : in_data <= 14'h0021; // 'd33
      10'd705  : in_data <= 14'h053b; // 'd1339
      10'd706  : in_data <= 14'h04d0; // 'd1232
      10'd707  : in_data <= 14'h0535; // 'd1333
      10'd708  : in_data <= 14'h01e2; // 'd482
      10'd709  : in_data <= 14'h0032; // 'd50
      10'd710  : in_data <= 14'h02cb; // 'd715
      10'd711  : in_data <= 14'h05a4; // 'd1444
      10'd712  : in_data <= 14'h0011; // 'd17
      10'd713  : in_data <= 14'h010e; // 'd270
      10'd714  : in_data <= 14'h045e; // 'd1118
      10'd715  : in_data <= 14'h05ee; // 'd1518
      10'd716  : in_data <= 14'h0354; // 'd852
      10'd717  : in_data <= 14'h051b; // 'd1307
      10'd718  : in_data <= 14'h0083; // 'd131
      10'd719  : in_data <= 14'h02fa; // 'd762
      10'd720  : in_data <= 14'h0440; // 'd1088
      10'd721  : in_data <= 14'h01cc; // 'd460
      10'd722  : in_data <= 14'h022f; // 'd559
      10'd723  : in_data <= 14'h0512; // 'd1298
      10'd724  : in_data <= 14'h04f7; // 'd1271
      10'd725  : in_data <= 14'h0395; // 'd917
      10'd726  : in_data <= 14'h032a; // 'd810
      10'd727  : in_data <= 14'h01c6; // 'd454
      10'd728  : in_data <= 14'h011e; // 'd286
      10'd729  : in_data <= 14'h0234; // 'd564
      10'd730  : in_data <= 14'h02b1; // 'd689
      10'd731  : in_data <= 14'h0093; // 'd147
      10'd732  : in_data <= 14'h0000; // 'd0
      10'd733  : in_data <= 14'h0066; // 'd102
      10'd734  : in_data <= 14'h0359; // 'd857
      10'd735  : in_data <= 14'h046d; // 'd1133
      10'd736  : in_data <= 14'h05af; // 'd1455
      10'd737  : in_data <= 14'h0069; // 'd105
      10'd738  : in_data <= 14'h05ad; // 'd1453
      10'd739  : in_data <= 14'h02dc; // 'd732
      10'd740  : in_data <= 14'h04a7; // 'd1191
      10'd741  : in_data <= 14'h010a; // 'd266
      10'd742  : in_data <= 14'h05ab; // 'd1451
      10'd743  : in_data <= 14'h0537; // 'd1335
      10'd744  : in_data <= 14'h00fa; // 'd250
      10'd745  : in_data <= 14'h05a0; // 'd1440
      10'd746  : in_data <= 14'h01ff; // 'd511
      10'd747  : in_data <= 14'h021d; // 'd541
      10'd748  : in_data <= 14'h0171; // 'd369
      10'd749  : in_data <= 14'h0117; // 'd279
      10'd750  : in_data <= 14'h00e3; // 'd227
      10'd751  : in_data <= 14'h02af; // 'd687
      10'd752  : in_data <= 14'h036b; // 'd875
      10'd753  : in_data <= 14'h04cd; // 'd1229
      10'd754  : in_data <= 14'h0347; // 'd839
      10'd755  : in_data <= 14'h0053; // 'd83
      10'd756  : in_data <= 14'h04d0; // 'd1232
      10'd757  : in_data <= 14'h02ba; // 'd698
      10'd758  : in_data <= 14'h04f4; // 'd1268
      10'd759  : in_data <= 14'h032f; // 'd815
      10'd760  : in_data <= 14'h006c; // 'd108
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      10'd0    : out_data_ref <= 8'h84;
      10'd1    : out_data_ref <= 8'hf3;
      10'd2    : out_data_ref <= 8'h27;
      10'd3    : out_data_ref <= 8'hd3;
      10'd4    : out_data_ref <= 8'h89;
      10'd5    : out_data_ref <= 8'h29;
      10'd6    : out_data_ref <= 8'h03;
      10'd7    : out_data_ref <= 8'h9e;
      10'd8    : out_data_ref <= 8'hf8;
      10'd9    : out_data_ref <= 8'h43;
      10'd10   : out_data_ref <= 8'h66;
      10'd11   : out_data_ref <= 8'hab;
      10'd12   : out_data_ref <= 8'h79;
      10'd13   : out_data_ref <= 8'h6a;
      10'd14   : out_data_ref <= 8'h96;
      10'd15   : out_data_ref <= 8'he6;
      10'd16   : out_data_ref <= 8'hcc;
      10'd17   : out_data_ref <= 8'h26;
      10'd18   : out_data_ref <= 8'h84;
      10'd19   : out_data_ref <= 8'h54;
      10'd20   : out_data_ref <= 8'hd5;
      10'd21   : out_data_ref <= 8'had;
      10'd22   : out_data_ref <= 8'h8d;
      10'd23   : out_data_ref <= 8'h05;
      10'd24   : out_data_ref <= 8'h41;
      10'd25   : out_data_ref <= 8'h0d;
      10'd26   : out_data_ref <= 8'h3e;
      10'd27   : out_data_ref <= 8'h96;
      10'd28   : out_data_ref <= 8'h9b;
      10'd29   : out_data_ref <= 8'h6d;
      10'd30   : out_data_ref <= 8'h22;
      10'd31   : out_data_ref <= 8'h8b;
      10'd32   : out_data_ref <= 8'h6c;
      10'd33   : out_data_ref <= 8'hed;
      10'd34   : out_data_ref <= 8'h2c;
      10'd35   : out_data_ref <= 8'hba;
      10'd36   : out_data_ref <= 8'hd7;
      10'd37   : out_data_ref <= 8'hba;
      10'd38   : out_data_ref <= 8'hb3;
      10'd39   : out_data_ref <= 8'hb4;
      10'd40   : out_data_ref <= 8'hb7;
      10'd41   : out_data_ref <= 8'hee;
      10'd42   : out_data_ref <= 8'h45;
      10'd43   : out_data_ref <= 8'h37;
      10'd44   : out_data_ref <= 8'h47;
      10'd45   : out_data_ref <= 8'hd3;
      10'd46   : out_data_ref <= 8'h33;
      10'd47   : out_data_ref <= 8'h1d;
      10'd48   : out_data_ref <= 8'h43;
      10'd49   : out_data_ref <= 8'hb2;
      10'd50   : out_data_ref <= 8'h1c;
      10'd51   : out_data_ref <= 8'hd2;
      10'd52   : out_data_ref <= 8'hec;
      10'd53   : out_data_ref <= 8'hc3;
      10'd54   : out_data_ref <= 8'hbf;
      10'd55   : out_data_ref <= 8'h55;
      10'd56   : out_data_ref <= 8'h7d;
      10'd57   : out_data_ref <= 8'h69;
      10'd58   : out_data_ref <= 8'h6e;
      10'd59   : out_data_ref <= 8'h81;
      10'd60   : out_data_ref <= 8'h77;
      10'd61   : out_data_ref <= 8'h3e;
      10'd62   : out_data_ref <= 8'he6;
      10'd63   : out_data_ref <= 8'h9f;
      10'd64   : out_data_ref <= 8'h68;
      10'd65   : out_data_ref <= 8'h7f;
      10'd66   : out_data_ref <= 8'he1;
      10'd67   : out_data_ref <= 8'hf6;
      10'd68   : out_data_ref <= 8'h1e;
      10'd69   : out_data_ref <= 8'h63;
      10'd70   : out_data_ref <= 8'h74;
      10'd71   : out_data_ref <= 8'h2a;
      10'd72   : out_data_ref <= 8'hf9;
      10'd73   : out_data_ref <= 8'h13;
      10'd74   : out_data_ref <= 8'ha3;
      10'd75   : out_data_ref <= 8'h54;
      10'd76   : out_data_ref <= 8'h18;
      10'd77   : out_data_ref <= 8'h57;
      10'd78   : out_data_ref <= 8'h54;
      10'd79   : out_data_ref <= 8'h67;
      10'd80   : out_data_ref <= 8'h11;
      10'd81   : out_data_ref <= 8'h84;
      10'd82   : out_data_ref <= 8'h09;
      10'd83   : out_data_ref <= 8'hd4;
      10'd84   : out_data_ref <= 8'hff;
      10'd85   : out_data_ref <= 8'hdb;
      10'd86   : out_data_ref <= 8'hba;
      10'd87   : out_data_ref <= 8'hc5;
      10'd88   : out_data_ref <= 8'hca;
      10'd89   : out_data_ref <= 8'h06;
      10'd90   : out_data_ref <= 8'h2d;
      10'd91   : out_data_ref <= 8'hff;
      10'd92   : out_data_ref <= 8'h3f;
      10'd93   : out_data_ref <= 8'h04;
      10'd94   : out_data_ref <= 8'hd7;
      10'd95   : out_data_ref <= 8'h61;
      10'd96   : out_data_ref <= 8'h54;
      10'd97   : out_data_ref <= 8'hd1;
      10'd98   : out_data_ref <= 8'h7e;
      10'd99   : out_data_ref <= 8'hc3;
      10'd100  : out_data_ref <= 8'h42;
      10'd101  : out_data_ref <= 8'h12;
      10'd102  : out_data_ref <= 8'hde;
      10'd103  : out_data_ref <= 8'hbf;
      10'd104  : out_data_ref <= 8'hca;
      10'd105  : out_data_ref <= 8'h96;
      10'd106  : out_data_ref <= 8'h7a;
      10'd107  : out_data_ref <= 8'h91;
      10'd108  : out_data_ref <= 8'he4;
      10'd109  : out_data_ref <= 8'h61;
      10'd110  : out_data_ref <= 8'hf7;
      10'd111  : out_data_ref <= 8'h37;
      10'd112  : out_data_ref <= 8'h86;
      10'd113  : out_data_ref <= 8'hd9;
      10'd114  : out_data_ref <= 8'h49;
      10'd115  : out_data_ref <= 8'hd6;
      10'd116  : out_data_ref <= 8'ha9;
      10'd117  : out_data_ref <= 8'h76;
      10'd118  : out_data_ref <= 8'h51;
      10'd119  : out_data_ref <= 8'h40;
      10'd120  : out_data_ref <= 8'hb9;
      10'd121  : out_data_ref <= 8'hdc;
      10'd122  : out_data_ref <= 8'h78;
      10'd123  : out_data_ref <= 8'h49;
      10'd124  : out_data_ref <= 8'h63;
      10'd125  : out_data_ref <= 8'h9a;
      10'd126  : out_data_ref <= 8'h48;
      10'd127  : out_data_ref <= 8'h70;
      10'd128  : out_data_ref <= 8'h58;
      10'd129  : out_data_ref <= 8'hf4;
      10'd130  : out_data_ref <= 8'h5d;
      10'd131  : out_data_ref <= 8'hda;
      10'd132  : out_data_ref <= 8'h91;
      10'd133  : out_data_ref <= 8'h95;
      10'd134  : out_data_ref <= 8'h76;
      10'd135  : out_data_ref <= 8'h09;
      10'd136  : out_data_ref <= 8'h0d;
      10'd137  : out_data_ref <= 8'h35;
      10'd138  : out_data_ref <= 8'he7;
      10'd139  : out_data_ref <= 8'h83;
      10'd140  : out_data_ref <= 8'h80;
      10'd141  : out_data_ref <= 8'h4b;
      10'd142  : out_data_ref <= 8'ha7;
      10'd143  : out_data_ref <= 8'hb8;
      10'd144  : out_data_ref <= 8'hb3;
      10'd145  : out_data_ref <= 8'h3b;
      10'd146  : out_data_ref <= 8'h5c;
      10'd147  : out_data_ref <= 8'h6a;
      10'd148  : out_data_ref <= 8'h8c;
      10'd149  : out_data_ref <= 8'h1e;
      10'd150  : out_data_ref <= 8'hbb;
      10'd151  : out_data_ref <= 8'h7c;
      10'd152  : out_data_ref <= 8'h39;
      10'd153  : out_data_ref <= 8'hf0;
      10'd154  : out_data_ref <= 8'h42;
      10'd155  : out_data_ref <= 8'h69;
      10'd156  : out_data_ref <= 8'h6c;
      10'd157  : out_data_ref <= 8'hf9;
      10'd158  : out_data_ref <= 8'hf2;
      10'd159  : out_data_ref <= 8'hb6;
      10'd160  : out_data_ref <= 8'h24;
      10'd161  : out_data_ref <= 8'hd2;
      10'd162  : out_data_ref <= 8'h6e;
      10'd163  : out_data_ref <= 8'ha5;
      10'd164  : out_data_ref <= 8'hd6;
      10'd165  : out_data_ref <= 8'hd1;
      10'd166  : out_data_ref <= 8'h01;
      10'd167  : out_data_ref <= 8'h48;
      10'd168  : out_data_ref <= 8'h9e;
      10'd169  : out_data_ref <= 8'h24;
      10'd170  : out_data_ref <= 8'h2c;
      10'd171  : out_data_ref <= 8'hc3;
      10'd172  : out_data_ref <= 8'h51;
      10'd173  : out_data_ref <= 8'h26;
      10'd174  : out_data_ref <= 8'hb5;
      10'd175  : out_data_ref <= 8'h73;
      10'd176  : out_data_ref <= 8'h92;
      10'd177  : out_data_ref <= 8'h8b;
      10'd178  : out_data_ref <= 8'h6b;
      10'd179  : out_data_ref <= 8'h8b;
      10'd180  : out_data_ref <= 8'hf9;
      10'd181  : out_data_ref <= 8'h94;
      10'd182  : out_data_ref <= 8'h52;
      10'd183  : out_data_ref <= 8'h69;
      10'd184  : out_data_ref <= 8'had;
      10'd185  : out_data_ref <= 8'h22;
      10'd186  : out_data_ref <= 8'he7;
      10'd187  : out_data_ref <= 8'hda;
      10'd188  : out_data_ref <= 8'h70;
      10'd189  : out_data_ref <= 8'hcc;
      10'd190  : out_data_ref <= 8'hb7;
      10'd191  : out_data_ref <= 8'hdc;
      10'd192  : out_data_ref <= 8'h37;
      10'd193  : out_data_ref <= 8'h4f;
      10'd194  : out_data_ref <= 8'h75;
      10'd195  : out_data_ref <= 8'h64;
      10'd196  : out_data_ref <= 8'h19;
      10'd197  : out_data_ref <= 8'h78;
      10'd198  : out_data_ref <= 8'hd5;
      10'd199  : out_data_ref <= 8'hf6;
      10'd200  : out_data_ref <= 8'hd5;
      10'd201  : out_data_ref <= 8'hf5;
      10'd202  : out_data_ref <= 8'h40;
      10'd203  : out_data_ref <= 8'ha1;
      10'd204  : out_data_ref <= 8'h16;
      10'd205  : out_data_ref <= 8'h9e;
      10'd206  : out_data_ref <= 8'hb0;
      10'd207  : out_data_ref <= 8'h98;
      10'd208  : out_data_ref <= 8'h57;
      10'd209  : out_data_ref <= 8'h0a;
      10'd210  : out_data_ref <= 8'h7c;
      10'd211  : out_data_ref <= 8'hfd;
      10'd212  : out_data_ref <= 8'h65;
      10'd213  : out_data_ref <= 8'hc9;
      10'd214  : out_data_ref <= 8'h25;
      10'd215  : out_data_ref <= 8'h7c;
      10'd216  : out_data_ref <= 8'h4c;
      10'd217  : out_data_ref <= 8'h19;
      10'd218  : out_data_ref <= 8'h6f;
      10'd219  : out_data_ref <= 8'h42;
      10'd220  : out_data_ref <= 8'hc6;
      10'd221  : out_data_ref <= 8'hda;
      10'd222  : out_data_ref <= 8'h4f;
      10'd223  : out_data_ref <= 8'h44;
      10'd224  : out_data_ref <= 8'h66;
      10'd225  : out_data_ref <= 8'hd8;
      10'd226  : out_data_ref <= 8'hf1;
      10'd227  : out_data_ref <= 8'h1a;
      10'd228  : out_data_ref <= 8'h17;
      10'd229  : out_data_ref <= 8'hc6;
      10'd230  : out_data_ref <= 8'ha7;
      10'd231  : out_data_ref <= 8'h5a;
      10'd232  : out_data_ref <= 8'h9b;
      10'd233  : out_data_ref <= 8'hdd;
      10'd234  : out_data_ref <= 8'h45;
      10'd235  : out_data_ref <= 8'hb5;
      10'd236  : out_data_ref <= 8'hac;
      10'd237  : out_data_ref <= 8'h77;
      10'd238  : out_data_ref <= 8'ha8;
      10'd239  : out_data_ref <= 8'h36;
      10'd240  : out_data_ref <= 8'h7b;
      10'd241  : out_data_ref <= 8'h00;
      10'd242  : out_data_ref <= 8'h5e;
      10'd243  : out_data_ref <= 8'hd2;
      10'd244  : out_data_ref <= 8'h21;
      10'd245  : out_data_ref <= 8'h41;
      10'd246  : out_data_ref <= 8'ha8;
      10'd247  : out_data_ref <= 8'h1b;
      10'd248  : out_data_ref <= 8'h99;
      10'd249  : out_data_ref <= 8'h5a;
      10'd250  : out_data_ref <= 8'h19;
      10'd251  : out_data_ref <= 8'he4;
      10'd252  : out_data_ref <= 8'hdc;
      10'd253  : out_data_ref <= 8'h9e;
      10'd254  : out_data_ref <= 8'h67;
      10'd255  : out_data_ref <= 8'h43;
      10'd256  : out_data_ref <= 8'hb4;
      10'd257  : out_data_ref <= 8'hb4;
      10'd258  : out_data_ref <= 8'h5e;
      10'd259  : out_data_ref <= 8'h03;
      10'd260  : out_data_ref <= 8'h29;
      10'd261  : out_data_ref <= 8'he7;
      10'd262  : out_data_ref <= 8'ha0;
      10'd263  : out_data_ref <= 8'h0d;
      10'd264  : out_data_ref <= 8'h3f;
      10'd265  : out_data_ref <= 8'hf9;
      10'd266  : out_data_ref <= 8'h0c;
      10'd267  : out_data_ref <= 8'h7a;
      10'd268  : out_data_ref <= 8'h91;
      10'd269  : out_data_ref <= 8'h7c;
      10'd270  : out_data_ref <= 8'hdc;
      10'd271  : out_data_ref <= 8'h9c;
      10'd272  : out_data_ref <= 8'ha7;
      10'd273  : out_data_ref <= 8'h5a;
      10'd274  : out_data_ref <= 8'h34;
      10'd275  : out_data_ref <= 8'hff;
      10'd276  : out_data_ref <= 8'hfd;
      10'd277  : out_data_ref <= 8'hd9;
      10'd278  : out_data_ref <= 8'ha3;
      10'd279  : out_data_ref <= 8'h21;
      10'd280  : out_data_ref <= 8'h75;
      10'd281  : out_data_ref <= 8'h1b;
      10'd282  : out_data_ref <= 8'h5c;
      10'd283  : out_data_ref <= 8'h8b;
      10'd284  : out_data_ref <= 8'h2a;
      10'd285  : out_data_ref <= 8'hb9;
      10'd286  : out_data_ref <= 8'he1;
      10'd287  : out_data_ref <= 8'hea;
      10'd288  : out_data_ref <= 8'h03;
      10'd289  : out_data_ref <= 8'h7c;
      10'd290  : out_data_ref <= 8'hf4;
      10'd291  : out_data_ref <= 8'h5c;
      10'd292  : out_data_ref <= 8'h04;
      10'd293  : out_data_ref <= 8'hb4;
      10'd294  : out_data_ref <= 8'h12;
      10'd295  : out_data_ref <= 8'ha9;
      10'd296  : out_data_ref <= 8'h7f;
      10'd297  : out_data_ref <= 8'h52;
      10'd298  : out_data_ref <= 8'he7;
      10'd299  : out_data_ref <= 8'hc6;
      10'd300  : out_data_ref <= 8'hd6;
      10'd301  : out_data_ref <= 8'h65;
      10'd302  : out_data_ref <= 8'h08;
      10'd303  : out_data_ref <= 8'h45;
      10'd304  : out_data_ref <= 8'h6d;
      10'd305  : out_data_ref <= 8'h91;
      10'd306  : out_data_ref <= 8'h17;
      10'd307  : out_data_ref <= 8'h96;
      10'd308  : out_data_ref <= 8'h12;
      10'd309  : out_data_ref <= 8'h57;
      10'd310  : out_data_ref <= 8'hb4;
      10'd311  : out_data_ref <= 8'hf5;
      10'd312  : out_data_ref <= 8'h0b;
      10'd313  : out_data_ref <= 8'hb9;
      10'd314  : out_data_ref <= 8'hf5;
      10'd315  : out_data_ref <= 8'h00;
      10'd316  : out_data_ref <= 8'hde;
      10'd317  : out_data_ref <= 8'h99;
      10'd318  : out_data_ref <= 8'hb6;
      10'd319  : out_data_ref <= 8'hf0;
      10'd320  : out_data_ref <= 8'h61;
      10'd321  : out_data_ref <= 8'hc3;
      10'd322  : out_data_ref <= 8'h77;
      10'd323  : out_data_ref <= 8'hd4;
      10'd324  : out_data_ref <= 8'h4f;
      10'd325  : out_data_ref <= 8'h49;
      10'd326  : out_data_ref <= 8'h5d;
      10'd327  : out_data_ref <= 8'h71;
      10'd328  : out_data_ref <= 8'h1a;
      10'd329  : out_data_ref <= 8'hb2;
      10'd330  : out_data_ref <= 8'hed;
      10'd331  : out_data_ref <= 8'h3e;
      10'd332  : out_data_ref <= 8'h88;
      10'd333  : out_data_ref <= 8'hcc;
      10'd334  : out_data_ref <= 8'hf1;
      10'd335  : out_data_ref <= 8'h4d;
      10'd336  : out_data_ref <= 8'hf1;
      10'd337  : out_data_ref <= 8'h0f;
      10'd338  : out_data_ref <= 8'h8c;
      10'd339  : out_data_ref <= 8'h60;
      10'd340  : out_data_ref <= 8'hbd;
      10'd341  : out_data_ref <= 8'h00;
      10'd342  : out_data_ref <= 8'he2;
      10'd343  : out_data_ref <= 8'h9c;
      10'd344  : out_data_ref <= 8'hd8;
      10'd345  : out_data_ref <= 8'h3a;
      10'd346  : out_data_ref <= 8'hd1;
      10'd347  : out_data_ref <= 8'h60;
      10'd348  : out_data_ref <= 8'hfa;
      10'd349  : out_data_ref <= 8'hef;
      10'd350  : out_data_ref <= 8'h29;
      10'd351  : out_data_ref <= 8'h84;
      10'd352  : out_data_ref <= 8'hfa;
      10'd353  : out_data_ref <= 8'hc7;
      10'd354  : out_data_ref <= 8'he8;
      10'd355  : out_data_ref <= 8'h97;
      10'd356  : out_data_ref <= 8'hcb;
      10'd357  : out_data_ref <= 8'hb8;
      10'd358  : out_data_ref <= 8'hcd;
      10'd359  : out_data_ref <= 8'ha1;
      10'd360  : out_data_ref <= 8'h44;
      10'd361  : out_data_ref <= 8'hd5;
      10'd362  : out_data_ref <= 8'h0e;
      10'd363  : out_data_ref <= 8'h4c;
      10'd364  : out_data_ref <= 8'h1a;
      10'd365  : out_data_ref <= 8'hd2;
      10'd366  : out_data_ref <= 8'h02;
      10'd367  : out_data_ref <= 8'h38;
      10'd368  : out_data_ref <= 8'ha2;
      10'd369  : out_data_ref <= 8'h61;
      10'd370  : out_data_ref <= 8'h75;
      10'd371  : out_data_ref <= 8'h98;
      10'd372  : out_data_ref <= 8'hda;
      10'd373  : out_data_ref <= 8'h6e;
      10'd374  : out_data_ref <= 8'hfe;
      10'd375  : out_data_ref <= 8'h78;
      10'd376  : out_data_ref <= 8'h6a;
      10'd377  : out_data_ref <= 8'ha8;
      10'd378  : out_data_ref <= 8'h2e;
      10'd379  : out_data_ref <= 8'h09;
      10'd380  : out_data_ref <= 8'h31;
      10'd381  : out_data_ref <= 8'hb0;
      10'd382  : out_data_ref <= 8'hb5;
      10'd383  : out_data_ref <= 8'hd1;
      10'd384  : out_data_ref <= 8'ha7;
      10'd385  : out_data_ref <= 8'hfa;
      10'd386  : out_data_ref <= 8'h02;
      10'd387  : out_data_ref <= 8'h4b;
      10'd388  : out_data_ref <= 8'h85;
      10'd389  : out_data_ref <= 8'h63;
      10'd390  : out_data_ref <= 8'h53;
      10'd391  : out_data_ref <= 8'haf;
      10'd392  : out_data_ref <= 8'hae;
      10'd393  : out_data_ref <= 8'hdb;
      10'd394  : out_data_ref <= 8'h0a;
      10'd395  : out_data_ref <= 8'h11;
      10'd396  : out_data_ref <= 8'h50;
      10'd397  : out_data_ref <= 8'ha4;
      10'd398  : out_data_ref <= 8'h2d;
      10'd399  : out_data_ref <= 8'ha1;
      10'd400  : out_data_ref <= 8'h82;
      10'd401  : out_data_ref <= 8'h35;
      10'd402  : out_data_ref <= 8'h3c;
      10'd403  : out_data_ref <= 8'he5;
      10'd404  : out_data_ref <= 8'ha0;
      10'd405  : out_data_ref <= 8'h04;
      10'd406  : out_data_ref <= 8'h03;
      10'd407  : out_data_ref <= 8'hbb;
      10'd408  : out_data_ref <= 8'h6b;
      10'd409  : out_data_ref <= 8'h7a;
      10'd410  : out_data_ref <= 8'h13;
      10'd411  : out_data_ref <= 8'hef;
      10'd412  : out_data_ref <= 8'hfc;
      10'd413  : out_data_ref <= 8'h14;
      10'd414  : out_data_ref <= 8'hb0;
      10'd415  : out_data_ref <= 8'hfd;
      10'd416  : out_data_ref <= 8'h97;
      10'd417  : out_data_ref <= 8'he1;
      10'd418  : out_data_ref <= 8'h11;
      10'd419  : out_data_ref <= 8'h73;
      10'd420  : out_data_ref <= 8'h02;
      10'd421  : out_data_ref <= 8'hed;
      10'd422  : out_data_ref <= 8'h8a;
      10'd423  : out_data_ref <= 8'h66;
      10'd424  : out_data_ref <= 8'hfa;
      10'd425  : out_data_ref <= 8'hae;
      10'd426  : out_data_ref <= 8'hd8;
      10'd427  : out_data_ref <= 8'h8b;
      10'd428  : out_data_ref <= 8'h43;
      10'd429  : out_data_ref <= 8'hb3;
      10'd430  : out_data_ref <= 8'h4c;
      10'd431  : out_data_ref <= 8'hfc;
      10'd432  : out_data_ref <= 8'h73;
      10'd433  : out_data_ref <= 8'hcb;
      10'd434  : out_data_ref <= 8'h33;
      10'd435  : out_data_ref <= 8'he4;
      10'd436  : out_data_ref <= 8'h9a;
      10'd437  : out_data_ref <= 8'h4c;
      10'd438  : out_data_ref <= 8'h34;
      10'd439  : out_data_ref <= 8'hd0;
      10'd440  : out_data_ref <= 8'hbf;
      10'd441  : out_data_ref <= 8'hde;
      10'd442  : out_data_ref <= 8'he2;
      10'd443  : out_data_ref <= 8'hfe;
      10'd444  : out_data_ref <= 8'had;
      10'd445  : out_data_ref <= 8'hc2;
      10'd446  : out_data_ref <= 8'hb4;
      10'd447  : out_data_ref <= 8'hc8;
      10'd448  : out_data_ref <= 8'hbb;
      10'd449  : out_data_ref <= 8'h1e;
      10'd450  : out_data_ref <= 8'hc4;
      10'd451  : out_data_ref <= 8'h12;
      10'd452  : out_data_ref <= 8'h15;
      10'd453  : out_data_ref <= 8'h58;
      10'd454  : out_data_ref <= 8'h6f;
      10'd455  : out_data_ref <= 8'hc6;
      10'd456  : out_data_ref <= 8'h65;
      10'd457  : out_data_ref <= 8'h50;
      10'd458  : out_data_ref <= 8'hd4;
      10'd459  : out_data_ref <= 8'h96;
      10'd460  : out_data_ref <= 8'h37;
      10'd461  : out_data_ref <= 8'h33;
      10'd462  : out_data_ref <= 8'h05;
      10'd463  : out_data_ref <= 8'hb9;
      10'd464  : out_data_ref <= 8'h9c;
      10'd465  : out_data_ref <= 8'hee;
      10'd466  : out_data_ref <= 8'h25;
      10'd467  : out_data_ref <= 8'h4e;
      10'd468  : out_data_ref <= 8'hac;
      10'd469  : out_data_ref <= 8'h71;
      10'd470  : out_data_ref <= 8'hd3;
      10'd471  : out_data_ref <= 8'hcd;
      10'd472  : out_data_ref <= 8'hac;
      10'd473  : out_data_ref <= 8'h68;
      10'd474  : out_data_ref <= 8'h9a;
      10'd475  : out_data_ref <= 8'h77;
      10'd476  : out_data_ref <= 8'h70;
      10'd477  : out_data_ref <= 8'h62;
      10'd478  : out_data_ref <= 8'hac;
      10'd479  : out_data_ref <= 8'hae;
      10'd480  : out_data_ref <= 8'h65;
      10'd481  : out_data_ref <= 8'hb0;
      10'd482  : out_data_ref <= 8'h31;
      10'd483  : out_data_ref <= 8'hb5;
      10'd484  : out_data_ref <= 8'ha1;
      10'd485  : out_data_ref <= 8'ha9;
      10'd486  : out_data_ref <= 8'h73;
      10'd487  : out_data_ref <= 8'h83;
      10'd488  : out_data_ref <= 8'h5b;
      10'd489  : out_data_ref <= 8'he6;
      10'd490  : out_data_ref <= 8'ha4;
      10'd491  : out_data_ref <= 8'hbb;
      10'd492  : out_data_ref <= 8'h06;
      10'd493  : out_data_ref <= 8'h1f;
      10'd494  : out_data_ref <= 8'h17;
      10'd495  : out_data_ref <= 8'h85;
      10'd496  : out_data_ref <= 8'h31;
      10'd497  : out_data_ref <= 8'hc4;
      10'd498  : out_data_ref <= 8'h5d;
      10'd499  : out_data_ref <= 8'he3;
      10'd500  : out_data_ref <= 8'hb3;
      10'd501  : out_data_ref <= 8'h3e;
      10'd502  : out_data_ref <= 8'h77;
      10'd503  : out_data_ref <= 8'h63;
      10'd504  : out_data_ref <= 8'hb4;
      10'd505  : out_data_ref <= 8'h83;
      10'd506  : out_data_ref <= 8'h62;
      10'd507  : out_data_ref <= 8'h18;
      10'd508  : out_data_ref <= 8'h21;
      10'd509  : out_data_ref <= 8'he0;
      10'd510  : out_data_ref <= 8'h37;
      10'd511  : out_data_ref <= 8'hfe;
      10'd512  : out_data_ref <= 8'h5e;
      10'd513  : out_data_ref <= 8'hf4;
      10'd514  : out_data_ref <= 8'h8f;
      10'd515  : out_data_ref <= 8'hd9;
      10'd516  : out_data_ref <= 8'h71;
      10'd517  : out_data_ref <= 8'hd8;
      10'd518  : out_data_ref <= 8'hd2;
      10'd519  : out_data_ref <= 8'hbe;
      10'd520  : out_data_ref <= 8'hfd;
      10'd521  : out_data_ref <= 8'ha6;
      10'd522  : out_data_ref <= 8'h32;
      10'd523  : out_data_ref <= 8'h50;
      10'd524  : out_data_ref <= 8'he9;
      10'd525  : out_data_ref <= 8'hb1;
      10'd526  : out_data_ref <= 8'h18;
      10'd527  : out_data_ref <= 8'h1d;
      10'd528  : out_data_ref <= 8'h8b;
      10'd529  : out_data_ref <= 8'h80;
      10'd530  : out_data_ref <= 8'h86;
      10'd531  : out_data_ref <= 8'hbe;
      10'd532  : out_data_ref <= 8'hd9;
      10'd533  : out_data_ref <= 8'hcd;
      10'd534  : out_data_ref <= 8'ha8;
      10'd535  : out_data_ref <= 8'hcd;
      10'd536  : out_data_ref <= 8'he6;
      10'd537  : out_data_ref <= 8'h64;
      10'd538  : out_data_ref <= 8'h4c;
      10'd539  : out_data_ref <= 8'hde;
      10'd540  : out_data_ref <= 8'h8e;
      10'd541  : out_data_ref <= 8'hbf;
      10'd542  : out_data_ref <= 8'h7c;
      10'd543  : out_data_ref <= 8'h1f;
      10'd544  : out_data_ref <= 8'h10;
      10'd545  : out_data_ref <= 8'h38;
      10'd546  : out_data_ref <= 8'haf;
      10'd547  : out_data_ref <= 8'he7;
      10'd548  : out_data_ref <= 8'h98;
      10'd549  : out_data_ref <= 8'ha2;
      10'd550  : out_data_ref <= 8'ha4;
      10'd551  : out_data_ref <= 8'hc4;
      10'd552  : out_data_ref <= 8'h92;
      10'd553  : out_data_ref <= 8'hb6;
      10'd554  : out_data_ref <= 8'h03;
      10'd555  : out_data_ref <= 8'hb7;
      10'd556  : out_data_ref <= 8'hf4;
      10'd557  : out_data_ref <= 8'hf8;
      10'd558  : out_data_ref <= 8'h80;
      10'd559  : out_data_ref <= 8'h5d;
      10'd560  : out_data_ref <= 8'h0f;
      10'd561  : out_data_ref <= 8'hdf;
      10'd562  : out_data_ref <= 8'h19;
      10'd563  : out_data_ref <= 8'hd8;
      10'd564  : out_data_ref <= 8'h27;
      10'd565  : out_data_ref <= 8'h48;
      10'd566  : out_data_ref <= 8'h88;
      10'd567  : out_data_ref <= 8'hce;
      10'd568  : out_data_ref <= 8'hbe;
      10'd569  : out_data_ref <= 8'hc3;
      10'd570  : out_data_ref <= 8'h04;
      10'd571  : out_data_ref <= 8'h3c;
      10'd572  : out_data_ref <= 8'hc9;
      10'd573  : out_data_ref <= 8'hac;
      10'd574  : out_data_ref <= 8'hf0;
      10'd575  : out_data_ref <= 8'h24;
      10'd576  : out_data_ref <= 8'hbd;
      10'd577  : out_data_ref <= 8'h30;
      10'd578  : out_data_ref <= 8'hd8;
      10'd579  : out_data_ref <= 8'hb0;
      10'd580  : out_data_ref <= 8'hd2;
      10'd581  : out_data_ref <= 8'h8d;
      10'd582  : out_data_ref <= 8'h31;
      10'd583  : out_data_ref <= 8'h19;
      10'd584  : out_data_ref <= 8'h85;
      10'd585  : out_data_ref <= 8'h93;
      10'd586  : out_data_ref <= 8'h01;
      10'd587  : out_data_ref <= 8'h10;
      10'd588  : out_data_ref <= 8'h38;
      10'd589  : out_data_ref <= 8'h65;
      10'd590  : out_data_ref <= 8'h98;
      10'd591  : out_data_ref <= 8'h77;
      10'd592  : out_data_ref <= 8'h5c;
      10'd593  : out_data_ref <= 8'hf8;
      10'd594  : out_data_ref <= 8'h4e;
      10'd595  : out_data_ref <= 8'h08;
      10'd596  : out_data_ref <= 8'h48;
      10'd597  : out_data_ref <= 8'hb1;
      10'd598  : out_data_ref <= 8'h1e;
      10'd599  : out_data_ref <= 8'h09;
      10'd600  : out_data_ref <= 8'h09;
      10'd601  : out_data_ref <= 8'h05;
      10'd602  : out_data_ref <= 8'ha6;
      10'd603  : out_data_ref <= 8'h5f;
      10'd604  : out_data_ref <= 8'h56;
      10'd605  : out_data_ref <= 8'h14;
      10'd606  : out_data_ref <= 8'h2f;
      10'd607  : out_data_ref <= 8'hc1;
      10'd608  : out_data_ref <= 8'h7d;
      10'd609  : out_data_ref <= 8'h25;
      10'd610  : out_data_ref <= 8'h73;
      10'd611  : out_data_ref <= 8'h53;
      10'd612  : out_data_ref <= 8'h6f;
      10'd613  : out_data_ref <= 8'hc5;
      10'd614  : out_data_ref <= 8'h1e;
      10'd615  : out_data_ref <= 8'h7d;
      10'd616  : out_data_ref <= 8'h5b;
      10'd617  : out_data_ref <= 8'h2e;
      10'd618  : out_data_ref <= 8'h0f;
      10'd619  : out_data_ref <= 8'hf7;
      10'd620  : out_data_ref <= 8'hb0;
      10'd621  : out_data_ref <= 8'h94;
      10'd622  : out_data_ref <= 8'h71;
      10'd623  : out_data_ref <= 8'h15;
      10'd624  : out_data_ref <= 8'h50;
      10'd625  : out_data_ref <= 8'h08;
      10'd626  : out_data_ref <= 8'h56;
      10'd627  : out_data_ref <= 8'h11;
      10'd628  : out_data_ref <= 8'h56;
      10'd629  : out_data_ref <= 8'hfb;
      10'd630  : out_data_ref <= 8'hae;
      10'd631  : out_data_ref <= 8'hc2;
      10'd632  : out_data_ref <= 8'h15;
      10'd633  : out_data_ref <= 8'h03;
      10'd634  : out_data_ref <= 8'h1e;
      10'd635  : out_data_ref <= 8'hd0;
      10'd636  : out_data_ref <= 8'hd8;
      10'd637  : out_data_ref <= 8'h44;
      10'd638  : out_data_ref <= 8'heb;
      10'd639  : out_data_ref <= 8'h14;
      10'd640  : out_data_ref <= 8'hd6;
      10'd641  : out_data_ref <= 8'hc6;
      10'd642  : out_data_ref <= 8'h09;
      10'd643  : out_data_ref <= 8'h17;
      10'd644  : out_data_ref <= 8'h33;
      10'd645  : out_data_ref <= 8'h55;
      10'd646  : out_data_ref <= 8'hff;
      10'd647  : out_data_ref <= 8'hf8;
      10'd648  : out_data_ref <= 8'hae;
      10'd649  : out_data_ref <= 8'h22;
      10'd650  : out_data_ref <= 8'hc6;
      10'd651  : out_data_ref <= 8'he5;
      10'd652  : out_data_ref <= 8'hbc;
      10'd653  : out_data_ref <= 8'hcd;
      10'd654  : out_data_ref <= 8'h19;
      10'd655  : out_data_ref <= 8'hb2;
      10'd656  : out_data_ref <= 8'h83;
      10'd657  : out_data_ref <= 8'h2e;
      10'd658  : out_data_ref <= 8'h5f;
      10'd659  : out_data_ref <= 8'hbe;
      10'd660  : out_data_ref <= 8'h62;
      10'd661  : out_data_ref <= 8'h5c;
      10'd662  : out_data_ref <= 8'h2c;
      10'd663  : out_data_ref <= 8'h0e;
      10'd664  : out_data_ref <= 8'h51;
      10'd665  : out_data_ref <= 8'h6e;
      10'd666  : out_data_ref <= 8'h13;
      10'd667  : out_data_ref <= 8'h69;
      10'd668  : out_data_ref <= 8'hd1;
      10'd669  : out_data_ref <= 8'hfc;
      10'd670  : out_data_ref <= 8'hf4;
      10'd671  : out_data_ref <= 8'h9a;
      10'd672  : out_data_ref <= 8'h5f;
      10'd673  : out_data_ref <= 8'hdb;
      10'd674  : out_data_ref <= 8'haf;
      10'd675  : out_data_ref <= 8'h8c;
      10'd676  : out_data_ref <= 8'hf5;
      10'd677  : out_data_ref <= 8'h72;
      10'd678  : out_data_ref <= 8'hf0;
      10'd679  : out_data_ref <= 8'h43;
      10'd680  : out_data_ref <= 8'h17;
      10'd681  : out_data_ref <= 8'hdb;
      10'd682  : out_data_ref <= 8'h8e;
      10'd683  : out_data_ref <= 8'hd7;
      10'd684  : out_data_ref <= 8'h0e;
      10'd685  : out_data_ref <= 8'he1;
      10'd686  : out_data_ref <= 8'h60;
      10'd687  : out_data_ref <= 8'h5b;
      10'd688  : out_data_ref <= 8'h96;
      10'd689  : out_data_ref <= 8'hd0;
      10'd690  : out_data_ref <= 8'h77;
      10'd691  : out_data_ref <= 8'hb4;
      10'd692  : out_data_ref <= 8'hf0;
      10'd693  : out_data_ref <= 8'h54;
      10'd694  : out_data_ref <= 8'hc7;
      10'd695  : out_data_ref <= 8'h2b;
      10'd696  : out_data_ref <= 8'h13;
      10'd697  : out_data_ref <= 8'h9f;
      10'd698  : out_data_ref <= 8'h5b;
      10'd699  : out_data_ref <= 8'hca;
      10'd700  : out_data_ref <= 8'ha5;
      10'd701  : out_data_ref <= 8'hbb;
      10'd702  : out_data_ref <= 8'h62;
      10'd703  : out_data_ref <= 8'h7e;
      10'd704  : out_data_ref <= 8'h39;
      10'd705  : out_data_ref <= 8'hbe;
      10'd706  : out_data_ref <= 8'h5b;
      10'd707  : out_data_ref <= 8'hcc;
      10'd708  : out_data_ref <= 8'h97;
      10'd709  : out_data_ref <= 8'haf;
      10'd710  : out_data_ref <= 8'h92;
      10'd711  : out_data_ref <= 8'h2c;
      10'd712  : out_data_ref <= 8'h5e;
      10'd713  : out_data_ref <= 8'h70;
      10'd714  : out_data_ref <= 8'h83;
      10'd715  : out_data_ref <= 8'h5b;
      10'd716  : out_data_ref <= 8'hd9;
      10'd717  : out_data_ref <= 8'h18;
      10'd718  : out_data_ref <= 8'h28;
      10'd719  : out_data_ref <= 8'h1b;
      10'd720  : out_data_ref <= 8'h95;
      10'd721  : out_data_ref <= 8'he5;
      10'd722  : out_data_ref <= 8'h57;
      10'd723  : out_data_ref <= 8'hfc;
      10'd724  : out_data_ref <= 8'h86;
      10'd725  : out_data_ref <= 8'ha4;
      10'd726  : out_data_ref <= 8'h3c;
      10'd727  : out_data_ref <= 8'h75;
      10'd728  : out_data_ref <= 8'h98;
      10'd729  : out_data_ref <= 8'h0a;
      10'd730  : out_data_ref <= 8'h0d;
      10'd731  : out_data_ref <= 8'h9f;
      10'd732  : out_data_ref <= 8'h0f;
      10'd733  : out_data_ref <= 8'h91;
      10'd734  : out_data_ref <= 8'h62;
      10'd735  : out_data_ref <= 8'hf2;
      10'd736  : out_data_ref <= 8'h30;
      10'd737  : out_data_ref <= 8'h01;
      10'd738  : out_data_ref <= 8'h4c;
      10'd739  : out_data_ref <= 8'hd8;
      10'd740  : out_data_ref <= 8'h67;
      10'd741  : out_data_ref <= 8'hdd;
      10'd742  : out_data_ref <= 8'h07;
      10'd743  : out_data_ref <= 8'hdb;
      10'd744  : out_data_ref <= 8'h23;
      10'd745  : out_data_ref <= 8'h26;
      10'd746  : out_data_ref <= 8'h09;
      10'd747  : out_data_ref <= 8'h34;
      10'd748  : out_data_ref <= 8'h54;
      10'd749  : out_data_ref <= 8'h6c;
      10'd750  : out_data_ref <= 8'h04;
      10'd751  : out_data_ref <= 8'h49;
      10'd752  : out_data_ref <= 8'h9d;
      10'd753  : out_data_ref <= 8'h6b;
      10'd754  : out_data_ref <= 8'h86;
      10'd755  : out_data_ref <= 8'h27;
      10'd756  : out_data_ref <= 8'hb8;
      10'd757  : out_data_ref <= 8'hd5;
      10'd758  : out_data_ref <= 8'hde;
      10'd759  : out_data_ref <= 8'hc7;
      10'd760  : out_data_ref <= 8'h3f;
      10'd761  : out_data_ref <= 8'ha4;
      10'd762  : out_data_ref <= 8'h53;
      10'd763  : out_data_ref <= 8'h27;
      10'd764  : out_data_ref <= 8'hf8;
      10'd765  : out_data_ref <= 8'h49;
      10'd766  : out_data_ref <= 8'h83;
      10'd767  : out_data_ref <= 8'h52;
      10'd768  : out_data_ref <= 8'h9b;
      10'd769  : out_data_ref <= 8'haf;
      10'd770  : out_data_ref <= 8'h3a;
      10'd771  : out_data_ref <= 8'ha1;
      10'd772  : out_data_ref <= 8'h0e;
      10'd773  : out_data_ref <= 8'h88;
      10'd774  : out_data_ref <= 8'h57;
      10'd775  : out_data_ref <= 8'h24;
      10'd776  : out_data_ref <= 8'hfe;
      10'd777  : out_data_ref <= 8'h76;
      10'd778  : out_data_ref <= 8'h05;
      10'd779  : out_data_ref <= 8'h50;
      10'd780  : out_data_ref <= 8'h99;
      10'd781  : out_data_ref <= 8'hd1;
      10'd782  : out_data_ref <= 8'h36;
      10'd783  : out_data_ref <= 8'hcc;
      10'd784  : out_data_ref <= 8'haa;
      10'd785  : out_data_ref <= 8'hcc;
      10'd786  : out_data_ref <= 8'h15;
      10'd787  : out_data_ref <= 8'h9b;
      10'd788  : out_data_ref <= 8'h4c;
      10'd789  : out_data_ref <= 8'he3;
      10'd790  : out_data_ref <= 8'h87;
      10'd791  : out_data_ref <= 8'h84;
      10'd792  : out_data_ref <= 8'h40;
      10'd793  : out_data_ref <= 8'h4c;
      10'd794  : out_data_ref <= 8'hc9;
      10'd795  : out_data_ref <= 8'hb0;
      10'd796  : out_data_ref <= 8'h47;
      10'd797  : out_data_ref <= 8'h23;
      10'd798  : out_data_ref <= 8'h91;
      10'd799  : out_data_ref <= 8'h0f;
      10'd800  : out_data_ref <= 8'h99;
      10'd801  : out_data_ref <= 8'h0a;
      10'd802  : out_data_ref <= 8'hf7;
      10'd803  : out_data_ref <= 8'h7c;
      10'd804  : out_data_ref <= 8'h64;
      10'd805  : out_data_ref <= 8'hd4;
      10'd806  : out_data_ref <= 8'h2a;
      10'd807  : out_data_ref <= 8'h29;
      10'd808  : out_data_ref <= 8'hd7;
      10'd809  : out_data_ref <= 8'h84;
      10'd810  : out_data_ref <= 8'hfc;
      10'd811  : out_data_ref <= 8'h89;
      10'd812  : out_data_ref <= 8'h79;
      10'd813  : out_data_ref <= 8'h55;
      10'd814  : out_data_ref <= 8'h75;
      10'd815  : out_data_ref <= 8'h8f;
      10'd816  : out_data_ref <= 8'h1d;
      10'd817  : out_data_ref <= 8'h2a;
      10'd818  : out_data_ref <= 8'h12;
      10'd819  : out_data_ref <= 8'hbb;
      10'd820  : out_data_ref <= 8'h7c;
      10'd821  : out_data_ref <= 8'h6f;
      10'd822  : out_data_ref <= 8'h6a;
      10'd823  : out_data_ref <= 8'h8e;
      10'd824  : out_data_ref <= 8'h5b;
      10'd825  : out_data_ref <= 8'h94;
      10'd826  : out_data_ref <= 8'hef;
      10'd827  : out_data_ref <= 8'ha7;
      10'd828  : out_data_ref <= 8'h40;
      10'd829  : out_data_ref <= 8'hf6;
      10'd830  : out_data_ref <= 8'h62;
      10'd831  : out_data_ref <= 8'hcf;
      10'd832  : out_data_ref <= 8'h0d;
      10'd833  : out_data_ref <= 8'ha2;
      10'd834  : out_data_ref <= 8'hd0;
      10'd835  : out_data_ref <= 8'h99;
      10'd836  : out_data_ref <= 8'hc6;
      10'd837  : out_data_ref <= 8'h1e;
      10'd838  : out_data_ref <= 8'he1;
      10'd839  : out_data_ref <= 8'hcc;
      10'd840  : out_data_ref <= 8'h6b;
      10'd841  : out_data_ref <= 8'h66;
      10'd842  : out_data_ref <= 8'h1a;
      10'd843  : out_data_ref <= 8'h64;
      10'd844  : out_data_ref <= 8'hf0;
      10'd845  : out_data_ref <= 8'h88;
      10'd846  : out_data_ref <= 8'h7b;
      10'd847  : out_data_ref <= 8'h80;
      10'd848  : out_data_ref <= 8'h5a;
      10'd849  : out_data_ref <= 8'hf5;
      10'd850  : out_data_ref <= 8'h3c;
      10'd851  : out_data_ref <= 8'h7b;
      10'd852  : out_data_ref <= 8'h64;
      10'd853  : out_data_ref <= 8'hc4;
      10'd854  : out_data_ref <= 8'h45;
      10'd855  : out_data_ref <= 8'h6d;
      10'd856  : out_data_ref <= 8'haf;
      10'd857  : out_data_ref <= 8'h22;
      10'd858  : out_data_ref <= 8'h85;
      10'd859  : out_data_ref <= 8'h82;
      10'd860  : out_data_ref <= 8'hc1;
      10'd861  : out_data_ref <= 8'hb2;
      10'd862  : out_data_ref <= 8'h21;
      10'd863  : out_data_ref <= 8'h2a;
      10'd864  : out_data_ref <= 8'h8f;
      10'd865  : out_data_ref <= 8'h71;
      10'd866  : out_data_ref <= 8'h8e;
      10'd867  : out_data_ref <= 8'h56;
      10'd868  : out_data_ref <= 8'hdf;
      10'd869  : out_data_ref <= 8'h6b;
      10'd870  : out_data_ref <= 8'h72;
      10'd871  : out_data_ref <= 8'hd7;
      10'd872  : out_data_ref <= 8'hef;
      10'd873  : out_data_ref <= 8'ha0;
      10'd874  : out_data_ref <= 8'hc5;
      10'd875  : out_data_ref <= 8'hd2;
      10'd876  : out_data_ref <= 8'h65;
      10'd877  : out_data_ref <= 8'h82;
      10'd878  : out_data_ref <= 8'hce;
      10'd879  : out_data_ref <= 8'h96;
      10'd880  : out_data_ref <= 8'hae;
      10'd881  : out_data_ref <= 8'hfc;
      10'd882  : out_data_ref <= 8'he1;
      10'd883  : out_data_ref <= 8'h3c;
      10'd884  : out_data_ref <= 8'hb2;
      10'd885  : out_data_ref <= 8'h83;
      10'd886  : out_data_ref <= 8'h0c;
      10'd887  : out_data_ref <= 8'h3f;
      10'd888  : out_data_ref <= 8'hb3;
      10'd889  : out_data_ref <= 8'h2e;
      10'd890  : out_data_ref <= 8'h51;
      10'd891  : out_data_ref <= 8'h15;
      10'd892  : out_data_ref <= 8'haa;
      10'd893  : out_data_ref <= 8'hcc;
      10'd894  : out_data_ref <= 8'h20;
      10'd895  : out_data_ref <= 8'hd3;
      10'd896  : out_data_ref <= 8'ha3;
      10'd897  : out_data_ref <= 8'h35;
      10'd898  : out_data_ref <= 8'hf7;
      10'd899  : out_data_ref <= 8'ha4;
      10'd900  : out_data_ref <= 8'hc1;
      10'd901  : out_data_ref <= 8'h2e;
      10'd902  : out_data_ref <= 8'h0c;
      10'd903  : out_data_ref <= 8'hd1;
      10'd904  : out_data_ref <= 8'hde;
      10'd905  : out_data_ref <= 8'h53;
      10'd906  : out_data_ref <= 8'h2d;
      10'd907  : out_data_ref <= 8'h8d;
      10'd908  : out_data_ref <= 8'h9d;
      10'd909  : out_data_ref <= 8'h42;
      10'd910  : out_data_ref <= 8'hd6;
      10'd911  : out_data_ref <= 8'h9b;
      10'd912  : out_data_ref <= 8'hc2;
      10'd913  : out_data_ref <= 8'hd0;
      10'd914  : out_data_ref <= 8'hbe;
      10'd915  : out_data_ref <= 8'h0a;
      10'd916  : out_data_ref <= 8'hc7;
      10'd917  : out_data_ref <= 8'hdf;
      10'd918  : out_data_ref <= 8'h3b;
      10'd919  : out_data_ref <= 8'h8f;
      10'd920  : out_data_ref <= 8'h41;
      10'd921  : out_data_ref <= 8'h6b;
      10'd922  : out_data_ref <= 8'h9a;
      10'd923  : out_data_ref <= 8'h53;
      10'd924  : out_data_ref <= 8'hdb;
      10'd925  : out_data_ref <= 8'h26;
      10'd926  : out_data_ref <= 8'h1c;
      10'd927  : out_data_ref <= 8'h47;
      10'd928  : out_data_ref <= 8'h27;
      10'd929  : out_data_ref <= 8'h27;
      10'd930  : out_data_ref <= 8'h25;
      10'd931  : out_data_ref <= 8'ha8;
      10'd932  : out_data_ref <= 8'ha8;
      10'd933  : out_data_ref <= 8'h82;
      10'd934  : out_data_ref <= 8'h98;
      10'd935  : out_data_ref <= 8'h67;
      10'd936  : out_data_ref <= 8'h83;
      10'd937  : out_data_ref <= 8'h51;
      10'd938  : out_data_ref <= 8'hb4;
      10'd939  : out_data_ref <= 8'h21;
      10'd940  : out_data_ref <= 8'h03;
      10'd941  : out_data_ref <= 8'h21;
      10'd942  : out_data_ref <= 8'h90;
      10'd943  : out_data_ref <= 8'h92;
      10'd944  : out_data_ref <= 8'h07;
      10'd945  : out_data_ref <= 8'h6b;
      10'd946  : out_data_ref <= 8'h6e;
      10'd947  : out_data_ref <= 8'hce;
      10'd948  : out_data_ref <= 8'h74;
      10'd949  : out_data_ref <= 8'h4d;
      10'd950  : out_data_ref <= 8'h99;
      10'd951  : out_data_ref <= 8'h33;
      10'd952  : out_data_ref <= 8'h88;
      10'd953  : out_data_ref <= 8'ha8;
      10'd954  : out_data_ref <= 8'hf2;
      10'd955  : out_data_ref <= 8'hc4;
      10'd956  : out_data_ref <= 8'h75;
      10'd957  : out_data_ref <= 8'h07;
      10'd958  : out_data_ref <= 8'h9c;
      10'd959  : out_data_ref <= 8'hb8;
      10'd960  : out_data_ref <= 8'hbc;
      10'd961  : out_data_ref <= 8'h4d;
      10'd962  : out_data_ref <= 8'hc4;
      10'd963  : out_data_ref <= 8'h92;
      10'd964  : out_data_ref <= 8'ha4;
      10'd965  : out_data_ref <= 8'h79;
      10'd966  : out_data_ref <= 8'h71;
      10'd967  : out_data_ref <= 8'h47;
      10'd968  : out_data_ref <= 8'hc0;
      10'd969  : out_data_ref <= 8'h1e;
      10'd970  : out_data_ref <= 8'ha3;
      10'd971  : out_data_ref <= 8'h50;
      10'd972  : out_data_ref <= 8'h82;
      10'd973  : out_data_ref <= 8'h25;
      10'd974  : out_data_ref <= 8'h82;
      10'd975  : out_data_ref <= 8'h6f;
      10'd976  : out_data_ref <= 8'h7a;
      10'd977  : out_data_ref <= 8'h3d;
      10'd978  : out_data_ref <= 8'h32;
      10'd979  : out_data_ref <= 8'hbf;
      10'd980  : out_data_ref <= 8'h50;
      10'd981  : out_data_ref <= 8'h2b;
      10'd982  : out_data_ref <= 8'h0f;
      10'd983  : out_data_ref <= 8'h45;
      10'd984  : out_data_ref <= 8'h52;
      10'd985  : out_data_ref <= 8'hf3;
      10'd986  : out_data_ref <= 8'h6f;
      10'd987  : out_data_ref <= 8'hc9;
      10'd988  : out_data_ref <= 8'hf6;
      10'd989  : out_data_ref <= 8'hfb;
      10'd990  : out_data_ref <= 8'h91;
      10'd991  : out_data_ref <= 8'he8;
      10'd992  : out_data_ref <= 8'h2d;
      10'd993  : out_data_ref <= 8'hb1;
      10'd994  : out_data_ref <= 8'h94;
      10'd995  : out_data_ref <= 8'h93;
      10'd996  : out_data_ref <= 8'h38;
      10'd997  : out_data_ref <= 8'hb4;
      10'd998  : out_data_ref <= 8'h54;
      10'd999  : out_data_ref <= 8'h36;
      10'd1000 : out_data_ref <= 8'hec;
      10'd1001 : out_data_ref <= 8'h0f;
      10'd1002 : out_data_ref <= 8'hf6;
      10'd1003 : out_data_ref <= 8'h3b;
      10'd1004 : out_data_ref <= 8'h53;
      10'd1005 : out_data_ref <= 8'hf9;
      10'd1006 : out_data_ref <= 8'h00;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
