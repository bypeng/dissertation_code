module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd761;
  localparam R_DEPTH = 'd10;
  localparam B_LEN = 'd1158;
  localparam B_DEPTH = 'd11;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [13: 0] in_data;
  input      [10: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 14'h10c8; // 'd4296
      10'd1    : in_data <= 14'h0472; // 'd1138
      10'd2    : in_data <= 14'h00b5; // 'd181
      10'd3    : in_data <= 14'h008c; // 'd140
      10'd4    : in_data <= 14'h0f34; // 'd3892
      10'd5    : in_data <= 14'h00e4; // 'd228
      10'd6    : in_data <= 14'h0d6c; // 'd3436
      10'd7    : in_data <= 14'h0866; // 'd2150
      10'd8    : in_data <= 14'h0ced; // 'd3309
      10'd9    : in_data <= 14'h0dd8; // 'd3544
      10'd10   : in_data <= 14'h0b60; // 'd2912
      10'd11   : in_data <= 14'h0629; // 'd1577
      10'd12   : in_data <= 14'h0fc1; // 'd4033
      10'd13   : in_data <= 14'h075d; // 'd1885
      10'd14   : in_data <= 14'h0520; // 'd1312
      10'd15   : in_data <= 14'h110b; // 'd4363
      10'd16   : in_data <= 14'h00fe; // 'd254
      10'd17   : in_data <= 14'h114f; // 'd4431
      10'd18   : in_data <= 14'h0ce0; // 'd3296
      10'd19   : in_data <= 14'h083e; // 'd2110
      10'd20   : in_data <= 14'h0053; // 'd83
      10'd21   : in_data <= 14'h0420; // 'd1056
      10'd22   : in_data <= 14'h115e; // 'd4446
      10'd23   : in_data <= 14'h11a8; // 'd4520
      10'd24   : in_data <= 14'h0557; // 'd1367
      10'd25   : in_data <= 14'h0535; // 'd1333
      10'd26   : in_data <= 14'h0920; // 'd2336
      10'd27   : in_data <= 14'h0a8e; // 'd2702
      10'd28   : in_data <= 14'h0804; // 'd2052
      10'd29   : in_data <= 14'h0463; // 'd1123
      10'd30   : in_data <= 14'h0c97; // 'd3223
      10'd31   : in_data <= 14'h0341; // 'd833
      10'd32   : in_data <= 14'h0e89; // 'd3721
      10'd33   : in_data <= 14'h104a; // 'd4170
      10'd34   : in_data <= 14'h0647; // 'd1607
      10'd35   : in_data <= 14'h03d5; // 'd981
      10'd36   : in_data <= 14'h064d; // 'd1613
      10'd37   : in_data <= 14'h055c; // 'd1372
      10'd38   : in_data <= 14'h0e37; // 'd3639
      10'd39   : in_data <= 14'h0890; // 'd2192
      10'd40   : in_data <= 14'h0f85; // 'd3973
      10'd41   : in_data <= 14'h054c; // 'd1356
      10'd42   : in_data <= 14'h0b33; // 'd2867
      10'd43   : in_data <= 14'h0466; // 'd1126
      10'd44   : in_data <= 14'h0795; // 'd1941
      10'd45   : in_data <= 14'h0a5d; // 'd2653
      10'd46   : in_data <= 14'h0081; // 'd129
      10'd47   : in_data <= 14'h0e75; // 'd3701
      10'd48   : in_data <= 14'h10f9; // 'd4345
      10'd49   : in_data <= 14'h0047; // 'd71
      10'd50   : in_data <= 14'h05bf; // 'd1471
      10'd51   : in_data <= 14'h10e7; // 'd4327
      10'd52   : in_data <= 14'h11c3; // 'd4547
      10'd53   : in_data <= 14'h08ee; // 'd2286
      10'd54   : in_data <= 14'h06f0; // 'd1776
      10'd55   : in_data <= 14'h0334; // 'd820
      10'd56   : in_data <= 14'h03e8; // 'd1000
      10'd57   : in_data <= 14'h0eb5; // 'd3765
      10'd58   : in_data <= 14'h0e36; // 'd3638
      10'd59   : in_data <= 14'h1000; // 'd4096
      10'd60   : in_data <= 14'h0aea; // 'd2794
      10'd61   : in_data <= 14'h026a; // 'd618
      10'd62   : in_data <= 14'h11e6; // 'd4582
      10'd63   : in_data <= 14'h0b48; // 'd2888
      10'd64   : in_data <= 14'h07ed; // 'd2029
      10'd65   : in_data <= 14'h0ee0; // 'd3808
      10'd66   : in_data <= 14'h00bf; // 'd191
      10'd67   : in_data <= 14'h06a8; // 'd1704
      10'd68   : in_data <= 14'h088b; // 'd2187
      10'd69   : in_data <= 14'h0de5; // 'd3557
      10'd70   : in_data <= 14'h0997; // 'd2455
      10'd71   : in_data <= 14'h03c5; // 'd965
      10'd72   : in_data <= 14'h100c; // 'd4108
      10'd73   : in_data <= 14'h0b5a; // 'd2906
      10'd74   : in_data <= 14'h0581; // 'd1409
      10'd75   : in_data <= 14'h098c; // 'd2444
      10'd76   : in_data <= 14'h00a0; // 'd160
      10'd77   : in_data <= 14'h096e; // 'd2414
      10'd78   : in_data <= 14'h0f31; // 'd3889
      10'd79   : in_data <= 14'h10cf; // 'd4303
      10'd80   : in_data <= 14'h0013; // 'd19
      10'd81   : in_data <= 14'h0dfc; // 'd3580
      10'd82   : in_data <= 14'h112c; // 'd4396
      10'd83   : in_data <= 14'h038e; // 'd910
      10'd84   : in_data <= 14'h0505; // 'd1285
      10'd85   : in_data <= 14'h0422; // 'd1058
      10'd86   : in_data <= 14'h0c36; // 'd3126
      10'd87   : in_data <= 14'h0d37; // 'd3383
      10'd88   : in_data <= 14'h0342; // 'd834
      10'd89   : in_data <= 14'h0901; // 'd2305
      10'd90   : in_data <= 14'h088b; // 'd2187
      10'd91   : in_data <= 14'h060d; // 'd1549
      10'd92   : in_data <= 14'h0575; // 'd1397
      10'd93   : in_data <= 14'h054d; // 'd1357
      10'd94   : in_data <= 14'h0674; // 'd1652
      10'd95   : in_data <= 14'h0a86; // 'd2694
      10'd96   : in_data <= 14'h118e; // 'd4494
      10'd97   : in_data <= 14'h1103; // 'd4355
      10'd98   : in_data <= 14'h090d; // 'd2317
      10'd99   : in_data <= 14'h0d50; // 'd3408
      10'd100  : in_data <= 14'h0ae4; // 'd2788
      10'd101  : in_data <= 14'h0e1e; // 'd3614
      10'd102  : in_data <= 14'h00b9; // 'd185
      10'd103  : in_data <= 14'h116f; // 'd4463
      10'd104  : in_data <= 14'h0ce9; // 'd3305
      10'd105  : in_data <= 14'h0a68; // 'd2664
      10'd106  : in_data <= 14'h009e; // 'd158
      10'd107  : in_data <= 14'h09e1; // 'd2529
      10'd108  : in_data <= 14'h08ab; // 'd2219
      10'd109  : in_data <= 14'h0c0e; // 'd3086
      10'd110  : in_data <= 14'h031d; // 'd797
      10'd111  : in_data <= 14'h04a8; // 'd1192
      10'd112  : in_data <= 14'h0e08; // 'd3592
      10'd113  : in_data <= 14'h044b; // 'd1099
      10'd114  : in_data <= 14'h0f19; // 'd3865
      10'd115  : in_data <= 14'h03ba; // 'd954
      10'd116  : in_data <= 14'h0894; // 'd2196
      10'd117  : in_data <= 14'h114f; // 'd4431
      10'd118  : in_data <= 14'h0f0b; // 'd3851
      10'd119  : in_data <= 14'h06bf; // 'd1727
      10'd120  : in_data <= 14'h080b; // 'd2059
      10'd121  : in_data <= 14'h0119; // 'd281
      10'd122  : in_data <= 14'h03f5; // 'd1013
      10'd123  : in_data <= 14'h0fdb; // 'd4059
      10'd124  : in_data <= 14'h0061; // 'd97
      10'd125  : in_data <= 14'h08d0; // 'd2256
      10'd126  : in_data <= 14'h04b4; // 'd1204
      10'd127  : in_data <= 14'h03a4; // 'd932
      10'd128  : in_data <= 14'h0330; // 'd816
      10'd129  : in_data <= 14'h112b; // 'd4395
      10'd130  : in_data <= 14'h104a; // 'd4170
      10'd131  : in_data <= 14'h0170; // 'd368
      10'd132  : in_data <= 14'h0247; // 'd583
      10'd133  : in_data <= 14'h051e; // 'd1310
      10'd134  : in_data <= 14'h0bc3; // 'd3011
      10'd135  : in_data <= 14'h03ea; // 'd1002
      10'd136  : in_data <= 14'h0937; // 'd2359
      10'd137  : in_data <= 14'h0579; // 'd1401
      10'd138  : in_data <= 14'h0f31; // 'd3889
      10'd139  : in_data <= 14'h0337; // 'd823
      10'd140  : in_data <= 14'h10ae; // 'd4270
      10'd141  : in_data <= 14'h04bb; // 'd1211
      10'd142  : in_data <= 14'h05a7; // 'd1447
      10'd143  : in_data <= 14'h01e9; // 'd489
      10'd144  : in_data <= 14'h0a6e; // 'd2670
      10'd145  : in_data <= 14'h10a7; // 'd4263
      10'd146  : in_data <= 14'h0e94; // 'd3732
      10'd147  : in_data <= 14'h0c52; // 'd3154
      10'd148  : in_data <= 14'h0976; // 'd2422
      10'd149  : in_data <= 14'h0eec; // 'd3820
      10'd150  : in_data <= 14'h08e5; // 'd2277
      10'd151  : in_data <= 14'h0383; // 'd899
      10'd152  : in_data <= 14'h0f2e; // 'd3886
      10'd153  : in_data <= 14'h0aa9; // 'd2729
      10'd154  : in_data <= 14'h0ce7; // 'd3303
      10'd155  : in_data <= 14'h0ccd; // 'd3277
      10'd156  : in_data <= 14'h1069; // 'd4201
      10'd157  : in_data <= 14'h0d02; // 'd3330
      10'd158  : in_data <= 14'h0e52; // 'd3666
      10'd159  : in_data <= 14'h00bb; // 'd187
      10'd160  : in_data <= 14'h0364; // 'd868
      10'd161  : in_data <= 14'h04a7; // 'd1191
      10'd162  : in_data <= 14'h0a81; // 'd2689
      10'd163  : in_data <= 14'h0984; // 'd2436
      10'd164  : in_data <= 14'h1006; // 'd4102
      10'd165  : in_data <= 14'h0fd0; // 'd4048
      10'd166  : in_data <= 14'h011e; // 'd286
      10'd167  : in_data <= 14'h06f1; // 'd1777
      10'd168  : in_data <= 14'h0b57; // 'd2903
      10'd169  : in_data <= 14'h0716; // 'd1814
      10'd170  : in_data <= 14'h03bb; // 'd955
      10'd171  : in_data <= 14'h0b7e; // 'd2942
      10'd172  : in_data <= 14'h0979; // 'd2425
      10'd173  : in_data <= 14'h11e3; // 'd4579
      10'd174  : in_data <= 14'h0f14; // 'd3860
      10'd175  : in_data <= 14'h03a4; // 'd932
      10'd176  : in_data <= 14'h1006; // 'd4102
      10'd177  : in_data <= 14'h0be3; // 'd3043
      10'd178  : in_data <= 14'h082f; // 'd2095
      10'd179  : in_data <= 14'h0175; // 'd373
      10'd180  : in_data <= 14'h08ef; // 'd2287
      10'd181  : in_data <= 14'h06ad; // 'd1709
      10'd182  : in_data <= 14'h079b; // 'd1947
      10'd183  : in_data <= 14'h001a; // 'd26
      10'd184  : in_data <= 14'h0f18; // 'd3864
      10'd185  : in_data <= 14'h0b5f; // 'd2911
      10'd186  : in_data <= 14'h0db0; // 'd3504
      10'd187  : in_data <= 14'h0c26; // 'd3110
      10'd188  : in_data <= 14'h0776; // 'd1910
      10'd189  : in_data <= 14'h0dbf; // 'd3519
      10'd190  : in_data <= 14'h0f0c; // 'd3852
      10'd191  : in_data <= 14'h0be0; // 'd3040
      10'd192  : in_data <= 14'h0cf6; // 'd3318
      10'd193  : in_data <= 14'h0609; // 'd1545
      10'd194  : in_data <= 14'h005e; // 'd94
      10'd195  : in_data <= 14'h0017; // 'd23
      10'd196  : in_data <= 14'h05ee; // 'd1518
      10'd197  : in_data <= 14'h0a74; // 'd2676
      10'd198  : in_data <= 14'h0adb; // 'd2779
      10'd199  : in_data <= 14'h0022; // 'd34
      10'd200  : in_data <= 14'h1178; // 'd4472
      10'd201  : in_data <= 14'h0370; // 'd880
      10'd202  : in_data <= 14'h01c9; // 'd457
      10'd203  : in_data <= 14'h033b; // 'd827
      10'd204  : in_data <= 14'h01f5; // 'd501
      10'd205  : in_data <= 14'h01bc; // 'd444
      10'd206  : in_data <= 14'h0d33; // 'd3379
      10'd207  : in_data <= 14'h0d05; // 'd3333
      10'd208  : in_data <= 14'h0d8b; // 'd3467
      10'd209  : in_data <= 14'h078b; // 'd1931
      10'd210  : in_data <= 14'h0c8b; // 'd3211
      10'd211  : in_data <= 14'h07d3; // 'd2003
      10'd212  : in_data <= 14'h0379; // 'd889
      10'd213  : in_data <= 14'h072c; // 'd1836
      10'd214  : in_data <= 14'h0739; // 'd1849
      10'd215  : in_data <= 14'h00f7; // 'd247
      10'd216  : in_data <= 14'h0935; // 'd2357
      10'd217  : in_data <= 14'h0fd7; // 'd4055
      10'd218  : in_data <= 14'h0033; // 'd51
      10'd219  : in_data <= 14'h1143; // 'd4419
      10'd220  : in_data <= 14'h0391; // 'd913
      10'd221  : in_data <= 14'h06c2; // 'd1730
      10'd222  : in_data <= 14'h0110; // 'd272
      10'd223  : in_data <= 14'h005c; // 'd92
      10'd224  : in_data <= 14'h058a; // 'd1418
      10'd225  : in_data <= 14'h0f8f; // 'd3983
      10'd226  : in_data <= 14'h005a; // 'd90
      10'd227  : in_data <= 14'h07b3; // 'd1971
      10'd228  : in_data <= 14'h028a; // 'd650
      10'd229  : in_data <= 14'h0569; // 'd1385
      10'd230  : in_data <= 14'h0118; // 'd280
      10'd231  : in_data <= 14'h0340; // 'd832
      10'd232  : in_data <= 14'h0fcf; // 'd4047
      10'd233  : in_data <= 14'h0ae6; // 'd2790
      10'd234  : in_data <= 14'h0cd1; // 'd3281
      10'd235  : in_data <= 14'h0ca3; // 'd3235
      10'd236  : in_data <= 14'h07ce; // 'd1998
      10'd237  : in_data <= 14'h0093; // 'd147
      10'd238  : in_data <= 14'h033c; // 'd828
      10'd239  : in_data <= 14'h0719; // 'd1817
      10'd240  : in_data <= 14'h006a; // 'd106
      10'd241  : in_data <= 14'h0ebc; // 'd3772
      10'd242  : in_data <= 14'h014b; // 'd331
      10'd243  : in_data <= 14'h0e9e; // 'd3742
      10'd244  : in_data <= 14'h0b7c; // 'd2940
      10'd245  : in_data <= 14'h090c; // 'd2316
      10'd246  : in_data <= 14'h008a; // 'd138
      10'd247  : in_data <= 14'h0881; // 'd2177
      10'd248  : in_data <= 14'h0cab; // 'd3243
      10'd249  : in_data <= 14'h08d3; // 'd2259
      10'd250  : in_data <= 14'h0cbb; // 'd3259
      10'd251  : in_data <= 14'h0499; // 'd1177
      10'd252  : in_data <= 14'h0e49; // 'd3657
      10'd253  : in_data <= 14'h0911; // 'd2321
      10'd254  : in_data <= 14'h0f86; // 'd3974
      10'd255  : in_data <= 14'h097c; // 'd2428
      10'd256  : in_data <= 14'h0ea6; // 'd3750
      10'd257  : in_data <= 14'h0349; // 'd841
      10'd258  : in_data <= 14'h06e3; // 'd1763
      10'd259  : in_data <= 14'h0643; // 'd1603
      10'd260  : in_data <= 14'h09e5; // 'd2533
      10'd261  : in_data <= 14'h0e74; // 'd3700
      10'd262  : in_data <= 14'h0312; // 'd786
      10'd263  : in_data <= 14'h0194; // 'd404
      10'd264  : in_data <= 14'h0477; // 'd1143
      10'd265  : in_data <= 14'h0575; // 'd1397
      10'd266  : in_data <= 14'h0883; // 'd2179
      10'd267  : in_data <= 14'h0fae; // 'd4014
      10'd268  : in_data <= 14'h02d8; // 'd728
      10'd269  : in_data <= 14'h00af; // 'd175
      10'd270  : in_data <= 14'h00cf; // 'd207
      10'd271  : in_data <= 14'h07fd; // 'd2045
      10'd272  : in_data <= 14'h0bb5; // 'd2997
      10'd273  : in_data <= 14'h05e9; // 'd1513
      10'd274  : in_data <= 14'h0a18; // 'd2584
      10'd275  : in_data <= 14'h0756; // 'd1878
      10'd276  : in_data <= 14'h04a6; // 'd1190
      10'd277  : in_data <= 14'h099a; // 'd2458
      10'd278  : in_data <= 14'h04cc; // 'd1228
      10'd279  : in_data <= 14'h0203; // 'd515
      10'd280  : in_data <= 14'h01a4; // 'd420
      10'd281  : in_data <= 14'h0679; // 'd1657
      10'd282  : in_data <= 14'h052a; // 'd1322
      10'd283  : in_data <= 14'h0ae3; // 'd2787
      10'd284  : in_data <= 14'h0e52; // 'd3666
      10'd285  : in_data <= 14'h0dc1; // 'd3521
      10'd286  : in_data <= 14'h10e5; // 'd4325
      10'd287  : in_data <= 14'h00cc; // 'd204
      10'd288  : in_data <= 14'h046f; // 'd1135
      10'd289  : in_data <= 14'h0289; // 'd649
      10'd290  : in_data <= 14'h0246; // 'd582
      10'd291  : in_data <= 14'h081a; // 'd2074
      10'd292  : in_data <= 14'h028e; // 'd654
      10'd293  : in_data <= 14'h0f56; // 'd3926
      10'd294  : in_data <= 14'h022f; // 'd559
      10'd295  : in_data <= 14'h005d; // 'd93
      10'd296  : in_data <= 14'h0e8b; // 'd3723
      10'd297  : in_data <= 14'h0cad; // 'd3245
      10'd298  : in_data <= 14'h09b2; // 'd2482
      10'd299  : in_data <= 14'h08f8; // 'd2296
      10'd300  : in_data <= 14'h0184; // 'd388
      10'd301  : in_data <= 14'h03b4; // 'd948
      10'd302  : in_data <= 14'h0fc5; // 'd4037
      10'd303  : in_data <= 14'h0870; // 'd2160
      10'd304  : in_data <= 14'h0eb4; // 'd3764
      10'd305  : in_data <= 14'h03b8; // 'd952
      10'd306  : in_data <= 14'h0b8d; // 'd2957
      10'd307  : in_data <= 14'h0f8f; // 'd3983
      10'd308  : in_data <= 14'h03f9; // 'd1017
      10'd309  : in_data <= 14'h068c; // 'd1676
      10'd310  : in_data <= 14'h0a3f; // 'd2623
      10'd311  : in_data <= 14'h0303; // 'd771
      10'd312  : in_data <= 14'h0f44; // 'd3908
      10'd313  : in_data <= 14'h1041; // 'd4161
      10'd314  : in_data <= 14'h076c; // 'd1900
      10'd315  : in_data <= 14'h0aac; // 'd2732
      10'd316  : in_data <= 14'h0cd9; // 'd3289
      10'd317  : in_data <= 14'h0fda; // 'd4058
      10'd318  : in_data <= 14'h026e; // 'd622
      10'd319  : in_data <= 14'h081f; // 'd2079
      10'd320  : in_data <= 14'h0f9e; // 'd3998
      10'd321  : in_data <= 14'h0038; // 'd56
      10'd322  : in_data <= 14'h08e3; // 'd2275
      10'd323  : in_data <= 14'h0bfa; // 'd3066
      10'd324  : in_data <= 14'h0837; // 'd2103
      10'd325  : in_data <= 14'h116c; // 'd4460
      10'd326  : in_data <= 14'h0329; // 'd809
      10'd327  : in_data <= 14'h1070; // 'd4208
      10'd328  : in_data <= 14'h0501; // 'd1281
      10'd329  : in_data <= 14'h0ecd; // 'd3789
      10'd330  : in_data <= 14'h01d5; // 'd469
      10'd331  : in_data <= 14'h0bb6; // 'd2998
      10'd332  : in_data <= 14'h0c6f; // 'd3183
      10'd333  : in_data <= 14'h044f; // 'd1103
      10'd334  : in_data <= 14'h07d1; // 'd2001
      10'd335  : in_data <= 14'h0904; // 'd2308
      10'd336  : in_data <= 14'h0db6; // 'd3510
      10'd337  : in_data <= 14'h0029; // 'd41
      10'd338  : in_data <= 14'h013e; // 'd318
      10'd339  : in_data <= 14'h0f31; // 'd3889
      10'd340  : in_data <= 14'h0829; // 'd2089
      10'd341  : in_data <= 14'h019b; // 'd411
      10'd342  : in_data <= 14'h03c8; // 'd968
      10'd343  : in_data <= 14'h0557; // 'd1367
      10'd344  : in_data <= 14'h1146; // 'd4422
      10'd345  : in_data <= 14'h0433; // 'd1075
      10'd346  : in_data <= 14'h0f77; // 'd3959
      10'd347  : in_data <= 14'h0fbc; // 'd4028
      10'd348  : in_data <= 14'h063d; // 'd1597
      10'd349  : in_data <= 14'h0226; // 'd550
      10'd350  : in_data <= 14'h0341; // 'd833
      10'd351  : in_data <= 14'h1047; // 'd4167
      10'd352  : in_data <= 14'h0c68; // 'd3176
      10'd353  : in_data <= 14'h0850; // 'd2128
      10'd354  : in_data <= 14'h09a4; // 'd2468
      10'd355  : in_data <= 14'h01c7; // 'd455
      10'd356  : in_data <= 14'h09d9; // 'd2521
      10'd357  : in_data <= 14'h09e9; // 'd2537
      10'd358  : in_data <= 14'h01d6; // 'd470
      10'd359  : in_data <= 14'h07c0; // 'd1984
      10'd360  : in_data <= 14'h0236; // 'd566
      10'd361  : in_data <= 14'h09f1; // 'd2545
      10'd362  : in_data <= 14'h0033; // 'd51
      10'd363  : in_data <= 14'h0347; // 'd839
      10'd364  : in_data <= 14'h10f0; // 'd4336
      10'd365  : in_data <= 14'h0132; // 'd306
      10'd366  : in_data <= 14'h08ed; // 'd2285
      10'd367  : in_data <= 14'h0d55; // 'd3413
      10'd368  : in_data <= 14'h04a2; // 'd1186
      10'd369  : in_data <= 14'h01f9; // 'd505
      10'd370  : in_data <= 14'h0dcc; // 'd3532
      10'd371  : in_data <= 14'h0302; // 'd770
      10'd372  : in_data <= 14'h1032; // 'd4146
      10'd373  : in_data <= 14'h0b5e; // 'd2910
      10'd374  : in_data <= 14'h0544; // 'd1348
      10'd375  : in_data <= 14'h03b5; // 'd949
      10'd376  : in_data <= 14'h050d; // 'd1293
      10'd377  : in_data <= 14'h0726; // 'd1830
      10'd378  : in_data <= 14'h0528; // 'd1320
      10'd379  : in_data <= 14'h0799; // 'd1945
      10'd380  : in_data <= 14'h0410; // 'd1040
      10'd381  : in_data <= 14'h0c3b; // 'd3131
      10'd382  : in_data <= 14'h006b; // 'd107
      10'd383  : in_data <= 14'h0e14; // 'd3604
      10'd384  : in_data <= 14'h0069; // 'd105
      10'd385  : in_data <= 14'h00db; // 'd219
      10'd386  : in_data <= 14'h0d15; // 'd3349
      10'd387  : in_data <= 14'h0261; // 'd609
      10'd388  : in_data <= 14'h0fa5; // 'd4005
      10'd389  : in_data <= 14'h0098; // 'd152
      10'd390  : in_data <= 14'h035d; // 'd861
      10'd391  : in_data <= 14'h1176; // 'd4470
      10'd392  : in_data <= 14'h0224; // 'd548
      10'd393  : in_data <= 14'h0d77; // 'd3447
      10'd394  : in_data <= 14'h0217; // 'd535
      10'd395  : in_data <= 14'h0418; // 'd1048
      10'd396  : in_data <= 14'h0660; // 'd1632
      10'd397  : in_data <= 14'h0db0; // 'd3504
      10'd398  : in_data <= 14'h05b8; // 'd1464
      10'd399  : in_data <= 14'h085d; // 'd2141
      10'd400  : in_data <= 14'h10e5; // 'd4325
      10'd401  : in_data <= 14'h1093; // 'd4243
      10'd402  : in_data <= 14'h03a5; // 'd933
      10'd403  : in_data <= 14'h0da3; // 'd3491
      10'd404  : in_data <= 14'h11e1; // 'd4577
      10'd405  : in_data <= 14'h11de; // 'd4574
      10'd406  : in_data <= 14'h0a3a; // 'd2618
      10'd407  : in_data <= 14'h106d; // 'd4205
      10'd408  : in_data <= 14'h0f4d; // 'd3917
      10'd409  : in_data <= 14'h078c; // 'd1932
      10'd410  : in_data <= 14'h03fb; // 'd1019
      10'd411  : in_data <= 14'h01bd; // 'd445
      10'd412  : in_data <= 14'h0ca2; // 'd3234
      10'd413  : in_data <= 14'h00bd; // 'd189
      10'd414  : in_data <= 14'h021a; // 'd538
      10'd415  : in_data <= 14'h05f0; // 'd1520
      10'd416  : in_data <= 14'h02a8; // 'd680
      10'd417  : in_data <= 14'h0ec8; // 'd3784
      10'd418  : in_data <= 14'h0fdd; // 'd4061
      10'd419  : in_data <= 14'h0818; // 'd2072
      10'd420  : in_data <= 14'h0242; // 'd578
      10'd421  : in_data <= 14'h024a; // 'd586
      10'd422  : in_data <= 14'h0804; // 'd2052
      10'd423  : in_data <= 14'h013e; // 'd318
      10'd424  : in_data <= 14'h0544; // 'd1348
      10'd425  : in_data <= 14'h04e6; // 'd1254
      10'd426  : in_data <= 14'h0607; // 'd1543
      10'd427  : in_data <= 14'h0a42; // 'd2626
      10'd428  : in_data <= 14'h07bb; // 'd1979
      10'd429  : in_data <= 14'h09e9; // 'd2537
      10'd430  : in_data <= 14'h01e8; // 'd488
      10'd431  : in_data <= 14'h0d0a; // 'd3338
      10'd432  : in_data <= 14'h0cb5; // 'd3253
      10'd433  : in_data <= 14'h06f0; // 'd1776
      10'd434  : in_data <= 14'h0693; // 'd1683
      10'd435  : in_data <= 14'h0479; // 'd1145
      10'd436  : in_data <= 14'h0d55; // 'd3413
      10'd437  : in_data <= 14'h0009; // 'd9
      10'd438  : in_data <= 14'h0878; // 'd2168
      10'd439  : in_data <= 14'h0f1e; // 'd3870
      10'd440  : in_data <= 14'h0177; // 'd375
      10'd441  : in_data <= 14'h06f4; // 'd1780
      10'd442  : in_data <= 14'h0c29; // 'd3113
      10'd443  : in_data <= 14'h03a7; // 'd935
      10'd444  : in_data <= 14'h0f9c; // 'd3996
      10'd445  : in_data <= 14'h0657; // 'd1623
      10'd446  : in_data <= 14'h0ba5; // 'd2981
      10'd447  : in_data <= 14'h06ef; // 'd1775
      10'd448  : in_data <= 14'h0194; // 'd404
      10'd449  : in_data <= 14'h11b4; // 'd4532
      10'd450  : in_data <= 14'h08ed; // 'd2285
      10'd451  : in_data <= 14'h1170; // 'd4464
      10'd452  : in_data <= 14'h03dd; // 'd989
      10'd453  : in_data <= 14'h053c; // 'd1340
      10'd454  : in_data <= 14'h0e91; // 'd3729
      10'd455  : in_data <= 14'h065d; // 'd1629
      10'd456  : in_data <= 14'h09a6; // 'd2470
      10'd457  : in_data <= 14'h0109; // 'd265
      10'd458  : in_data <= 14'h03f1; // 'd1009
      10'd459  : in_data <= 14'h0eff; // 'd3839
      10'd460  : in_data <= 14'h09a6; // 'd2470
      10'd461  : in_data <= 14'h118d; // 'd4493
      10'd462  : in_data <= 14'h0c51; // 'd3153
      10'd463  : in_data <= 14'h0f1d; // 'd3869
      10'd464  : in_data <= 14'h09b6; // 'd2486
      10'd465  : in_data <= 14'h0aac; // 'd2732
      10'd466  : in_data <= 14'h0ee9; // 'd3817
      10'd467  : in_data <= 14'h0e46; // 'd3654
      10'd468  : in_data <= 14'h113c; // 'd4412
      10'd469  : in_data <= 14'h0a24; // 'd2596
      10'd470  : in_data <= 14'h0fb4; // 'd4020
      10'd471  : in_data <= 14'h06b1; // 'd1713
      10'd472  : in_data <= 14'h06db; // 'd1755
      10'd473  : in_data <= 14'h0054; // 'd84
      10'd474  : in_data <= 14'h0467; // 'd1127
      10'd475  : in_data <= 14'h06cf; // 'd1743
      10'd476  : in_data <= 14'h1104; // 'd4356
      10'd477  : in_data <= 14'h09a7; // 'd2471
      10'd478  : in_data <= 14'h0b57; // 'd2903
      10'd479  : in_data <= 14'h05d5; // 'd1493
      10'd480  : in_data <= 14'h0e9a; // 'd3738
      10'd481  : in_data <= 14'h08ef; // 'd2287
      10'd482  : in_data <= 14'h01d8; // 'd472
      10'd483  : in_data <= 14'h0969; // 'd2409
      10'd484  : in_data <= 14'h0705; // 'd1797
      10'd485  : in_data <= 14'h05eb; // 'd1515
      10'd486  : in_data <= 14'h08ec; // 'd2284
      10'd487  : in_data <= 14'h0be6; // 'd3046
      10'd488  : in_data <= 14'h05f3; // 'd1523
      10'd489  : in_data <= 14'h0d4c; // 'd3404
      10'd490  : in_data <= 14'h0eb3; // 'd3763
      10'd491  : in_data <= 14'h0ae2; // 'd2786
      10'd492  : in_data <= 14'h0e63; // 'd3683
      10'd493  : in_data <= 14'h00d9; // 'd217
      10'd494  : in_data <= 14'h0a18; // 'd2584
      10'd495  : in_data <= 14'h02dd; // 'd733
      10'd496  : in_data <= 14'h0f38; // 'd3896
      10'd497  : in_data <= 14'h0301; // 'd769
      10'd498  : in_data <= 14'h1128; // 'd4392
      10'd499  : in_data <= 14'h088a; // 'd2186
      10'd500  : in_data <= 14'h09ce; // 'd2510
      10'd501  : in_data <= 14'h0fbb; // 'd4027
      10'd502  : in_data <= 14'h054a; // 'd1354
      10'd503  : in_data <= 14'h0dd1; // 'd3537
      10'd504  : in_data <= 14'h04eb; // 'd1259
      10'd505  : in_data <= 14'h0a99; // 'd2713
      10'd506  : in_data <= 14'h0d09; // 'd3337
      10'd507  : in_data <= 14'h06e0; // 'd1760
      10'd508  : in_data <= 14'h017c; // 'd380
      10'd509  : in_data <= 14'h0297; // 'd663
      10'd510  : in_data <= 14'h1172; // 'd4466
      10'd511  : in_data <= 14'h08ce; // 'd2254
      10'd512  : in_data <= 14'h0f28; // 'd3880
      10'd513  : in_data <= 14'h1083; // 'd4227
      10'd514  : in_data <= 14'h02dc; // 'd732
      10'd515  : in_data <= 14'h074b; // 'd1867
      10'd516  : in_data <= 14'h0d36; // 'd3382
      10'd517  : in_data <= 14'h0ded; // 'd3565
      10'd518  : in_data <= 14'h0991; // 'd2449
      10'd519  : in_data <= 14'h0535; // 'd1333
      10'd520  : in_data <= 14'h058f; // 'd1423
      10'd521  : in_data <= 14'h1065; // 'd4197
      10'd522  : in_data <= 14'h0817; // 'd2071
      10'd523  : in_data <= 14'h07aa; // 'd1962
      10'd524  : in_data <= 14'h0004; // 'd4
      10'd525  : in_data <= 14'h0c02; // 'd3074
      10'd526  : in_data <= 14'h0e3b; // 'd3643
      10'd527  : in_data <= 14'h0b6b; // 'd2923
      10'd528  : in_data <= 14'h10a9; // 'd4265
      10'd529  : in_data <= 14'h09d0; // 'd2512
      10'd530  : in_data <= 14'h0c03; // 'd3075
      10'd531  : in_data <= 14'h0b85; // 'd2949
      10'd532  : in_data <= 14'h0b05; // 'd2821
      10'd533  : in_data <= 14'h0fba; // 'd4026
      10'd534  : in_data <= 14'h102d; // 'd4141
      10'd535  : in_data <= 14'h0b9a; // 'd2970
      10'd536  : in_data <= 14'h066c; // 'd1644
      10'd537  : in_data <= 14'h04b2; // 'd1202
      10'd538  : in_data <= 14'h0c90; // 'd3216
      10'd539  : in_data <= 14'h08af; // 'd2223
      10'd540  : in_data <= 14'h0f4e; // 'd3918
      10'd541  : in_data <= 14'h0abf; // 'd2751
      10'd542  : in_data <= 14'h0350; // 'd848
      10'd543  : in_data <= 14'h0f89; // 'd3977
      10'd544  : in_data <= 14'h100e; // 'd4110
      10'd545  : in_data <= 14'h0d80; // 'd3456
      10'd546  : in_data <= 14'h0a59; // 'd2649
      10'd547  : in_data <= 14'h0e17; // 'd3607
      10'd548  : in_data <= 14'h07e1; // 'd2017
      10'd549  : in_data <= 14'h0206; // 'd518
      10'd550  : in_data <= 14'h085d; // 'd2141
      10'd551  : in_data <= 14'h0901; // 'd2305
      10'd552  : in_data <= 14'h092a; // 'd2346
      10'd553  : in_data <= 14'h05b0; // 'd1456
      10'd554  : in_data <= 14'h0783; // 'd1923
      10'd555  : in_data <= 14'h0e10; // 'd3600
      10'd556  : in_data <= 14'h0b6a; // 'd2922
      10'd557  : in_data <= 14'h0883; // 'd2179
      10'd558  : in_data <= 14'h0191; // 'd401
      10'd559  : in_data <= 14'h0e3e; // 'd3646
      10'd560  : in_data <= 14'h11aa; // 'd4522
      10'd561  : in_data <= 14'h0e11; // 'd3601
      10'd562  : in_data <= 14'h05f8; // 'd1528
      10'd563  : in_data <= 14'h0f7a; // 'd3962
      10'd564  : in_data <= 14'h084f; // 'd2127
      10'd565  : in_data <= 14'h076c; // 'd1900
      10'd566  : in_data <= 14'h01cf; // 'd463
      10'd567  : in_data <= 14'h0634; // 'd1588
      10'd568  : in_data <= 14'h0428; // 'd1064
      10'd569  : in_data <= 14'h0911; // 'd2321
      10'd570  : in_data <= 14'h0c2d; // 'd3117
      10'd571  : in_data <= 14'h02eb; // 'd747
      10'd572  : in_data <= 14'h06f8; // 'd1784
      10'd573  : in_data <= 14'h0286; // 'd646
      10'd574  : in_data <= 14'h0a29; // 'd2601
      10'd575  : in_data <= 14'h0fe8; // 'd4072
      10'd576  : in_data <= 14'h0ec2; // 'd3778
      10'd577  : in_data <= 14'h0391; // 'd913
      10'd578  : in_data <= 14'h0c23; // 'd3107
      10'd579  : in_data <= 14'h0d63; // 'd3427
      10'd580  : in_data <= 14'h0e4d; // 'd3661
      10'd581  : in_data <= 14'h0349; // 'd841
      10'd582  : in_data <= 14'h101e; // 'd4126
      10'd583  : in_data <= 14'h0885; // 'd2181
      10'd584  : in_data <= 14'h0298; // 'd664
      10'd585  : in_data <= 14'h0c0a; // 'd3082
      10'd586  : in_data <= 14'h0ddc; // 'd3548
      10'd587  : in_data <= 14'h0077; // 'd119
      10'd588  : in_data <= 14'h0340; // 'd832
      10'd589  : in_data <= 14'h0494; // 'd1172
      10'd590  : in_data <= 14'h0420; // 'd1056
      10'd591  : in_data <= 14'h0543; // 'd1347
      10'd592  : in_data <= 14'h102d; // 'd4141
      10'd593  : in_data <= 14'h093c; // 'd2364
      10'd594  : in_data <= 14'h0668; // 'd1640
      10'd595  : in_data <= 14'h0b11; // 'd2833
      10'd596  : in_data <= 14'h08d2; // 'd2258
      10'd597  : in_data <= 14'h10cb; // 'd4299
      10'd598  : in_data <= 14'h0d6c; // 'd3436
      10'd599  : in_data <= 14'h0785; // 'd1925
      10'd600  : in_data <= 14'h0062; // 'd98
      10'd601  : in_data <= 14'h0107; // 'd263
      10'd602  : in_data <= 14'h063c; // 'd1596
      10'd603  : in_data <= 14'h0fe7; // 'd4071
      10'd604  : in_data <= 14'h070a; // 'd1802
      10'd605  : in_data <= 14'h0621; // 'd1569
      10'd606  : in_data <= 14'h0746; // 'd1862
      10'd607  : in_data <= 14'h1050; // 'd4176
      10'd608  : in_data <= 14'h081c; // 'd2076
      10'd609  : in_data <= 14'h0c09; // 'd3081
      10'd610  : in_data <= 14'h107d; // 'd4221
      10'd611  : in_data <= 14'h0ce0; // 'd3296
      10'd612  : in_data <= 14'h1114; // 'd4372
      10'd613  : in_data <= 14'h05a2; // 'd1442
      10'd614  : in_data <= 14'h11b4; // 'd4532
      10'd615  : in_data <= 14'h072f; // 'd1839
      10'd616  : in_data <= 14'h03e4; // 'd996
      10'd617  : in_data <= 14'h096b; // 'd2411
      10'd618  : in_data <= 14'h1127; // 'd4391
      10'd619  : in_data <= 14'h10fa; // 'd4346
      10'd620  : in_data <= 14'h071b; // 'd1819
      10'd621  : in_data <= 14'h08bf; // 'd2239
      10'd622  : in_data <= 14'h0bda; // 'd3034
      10'd623  : in_data <= 14'h0050; // 'd80
      10'd624  : in_data <= 14'h0fa8; // 'd4008
      10'd625  : in_data <= 14'h0c23; // 'd3107
      10'd626  : in_data <= 14'h10f8; // 'd4344
      10'd627  : in_data <= 14'h062c; // 'd1580
      10'd628  : in_data <= 14'h02d0; // 'd720
      10'd629  : in_data <= 14'h0678; // 'd1656
      10'd630  : in_data <= 14'h0029; // 'd41
      10'd631  : in_data <= 14'h0cc5; // 'd3269
      10'd632  : in_data <= 14'h1078; // 'd4216
      10'd633  : in_data <= 14'h0d86; // 'd3462
      10'd634  : in_data <= 14'h095d; // 'd2397
      10'd635  : in_data <= 14'h09fd; // 'd2557
      10'd636  : in_data <= 14'h0873; // 'd2163
      10'd637  : in_data <= 14'h11a4; // 'd4516
      10'd638  : in_data <= 14'h1018; // 'd4120
      10'd639  : in_data <= 14'h040b; // 'd1035
      10'd640  : in_data <= 14'h0f5d; // 'd3933
      10'd641  : in_data <= 14'h109b; // 'd4251
      10'd642  : in_data <= 14'h10dc; // 'd4316
      10'd643  : in_data <= 14'h066c; // 'd1644
      10'd644  : in_data <= 14'h04d4; // 'd1236
      10'd645  : in_data <= 14'h10fc; // 'd4348
      10'd646  : in_data <= 14'h0ff8; // 'd4088
      10'd647  : in_data <= 14'h054d; // 'd1357
      10'd648  : in_data <= 14'h0aec; // 'd2796
      10'd649  : in_data <= 14'h024d; // 'd589
      10'd650  : in_data <= 14'h08bb; // 'd2235
      10'd651  : in_data <= 14'h00ca; // 'd202
      10'd652  : in_data <= 14'h0b9f; // 'd2975
      10'd653  : in_data <= 14'h08c7; // 'd2247
      10'd654  : in_data <= 14'h0669; // 'd1641
      10'd655  : in_data <= 14'h1065; // 'd4197
      10'd656  : in_data <= 14'h0c7d; // 'd3197
      10'd657  : in_data <= 14'h04de; // 'd1246
      10'd658  : in_data <= 14'h1088; // 'd4232
      10'd659  : in_data <= 14'h07fa; // 'd2042
      10'd660  : in_data <= 14'h0225; // 'd549
      10'd661  : in_data <= 14'h1033; // 'd4147
      10'd662  : in_data <= 14'h0c2d; // 'd3117
      10'd663  : in_data <= 14'h0ebd; // 'd3773
      10'd664  : in_data <= 14'h0692; // 'd1682
      10'd665  : in_data <= 14'h0399; // 'd921
      10'd666  : in_data <= 14'h08a5; // 'd2213
      10'd667  : in_data <= 14'h054d; // 'd1357
      10'd668  : in_data <= 14'h109c; // 'd4252
      10'd669  : in_data <= 14'h05ec; // 'd1516
      10'd670  : in_data <= 14'h0d70; // 'd3440
      10'd671  : in_data <= 14'h02ce; // 'd718
      10'd672  : in_data <= 14'h0eb9; // 'd3769
      10'd673  : in_data <= 14'h0ccd; // 'd3277
      10'd674  : in_data <= 14'h104e; // 'd4174
      10'd675  : in_data <= 14'h01c4; // 'd452
      10'd676  : in_data <= 14'h0c33; // 'd3123
      10'd677  : in_data <= 14'h0a6a; // 'd2666
      10'd678  : in_data <= 14'h0318; // 'd792
      10'd679  : in_data <= 14'h0e76; // 'd3702
      10'd680  : in_data <= 14'h0bcf; // 'd3023
      10'd681  : in_data <= 14'h045e; // 'd1118
      10'd682  : in_data <= 14'h0695; // 'd1685
      10'd683  : in_data <= 14'h097b; // 'd2427
      10'd684  : in_data <= 14'h0577; // 'd1399
      10'd685  : in_data <= 14'h0090; // 'd144
      10'd686  : in_data <= 14'h0670; // 'd1648
      10'd687  : in_data <= 14'h11b5; // 'd4533
      10'd688  : in_data <= 14'h033b; // 'd827
      10'd689  : in_data <= 14'h0b55; // 'd2901
      10'd690  : in_data <= 14'h0671; // 'd1649
      10'd691  : in_data <= 14'h0910; // 'd2320
      10'd692  : in_data <= 14'h0245; // 'd581
      10'd693  : in_data <= 14'h10ea; // 'd4330
      10'd694  : in_data <= 14'h01d5; // 'd469
      10'd695  : in_data <= 14'h0a8d; // 'd2701
      10'd696  : in_data <= 14'h0ac8; // 'd2760
      10'd697  : in_data <= 14'h0ab3; // 'd2739
      10'd698  : in_data <= 14'h0877; // 'd2167
      10'd699  : in_data <= 14'h0409; // 'd1033
      10'd700  : in_data <= 14'h0b94; // 'd2964
      10'd701  : in_data <= 14'h1054; // 'd4180
      10'd702  : in_data <= 14'h07bf; // 'd1983
      10'd703  : in_data <= 14'h11d5; // 'd4565
      10'd704  : in_data <= 14'h08d6; // 'd2262
      10'd705  : in_data <= 14'h0a26; // 'd2598
      10'd706  : in_data <= 14'h0b59; // 'd2905
      10'd707  : in_data <= 14'h052f; // 'd1327
      10'd708  : in_data <= 14'h0f42; // 'd3906
      10'd709  : in_data <= 14'h0fe7; // 'd4071
      10'd710  : in_data <= 14'h0ca2; // 'd3234
      10'd711  : in_data <= 14'h0b0e; // 'd2830
      10'd712  : in_data <= 14'h0a94; // 'd2708
      10'd713  : in_data <= 14'h0f54; // 'd3924
      10'd714  : in_data <= 14'h0591; // 'd1425
      10'd715  : in_data <= 14'h0f66; // 'd3942
      10'd716  : in_data <= 14'h03ad; // 'd941
      10'd717  : in_data <= 14'h0cbe; // 'd3262
      10'd718  : in_data <= 14'h101d; // 'd4125
      10'd719  : in_data <= 14'h0bc1; // 'd3009
      10'd720  : in_data <= 14'h040f; // 'd1039
      10'd721  : in_data <= 14'h0069; // 'd105
      10'd722  : in_data <= 14'h03ec; // 'd1004
      10'd723  : in_data <= 14'h0022; // 'd34
      10'd724  : in_data <= 14'h05a4; // 'd1444
      10'd725  : in_data <= 14'h0380; // 'd896
      10'd726  : in_data <= 14'h0ebd; // 'd3773
      10'd727  : in_data <= 14'h0e0a; // 'd3594
      10'd728  : in_data <= 14'h0c31; // 'd3121
      10'd729  : in_data <= 14'h073c; // 'd1852
      10'd730  : in_data <= 14'h0076; // 'd118
      10'd731  : in_data <= 14'h0b5e; // 'd2910
      10'd732  : in_data <= 14'h0b57; // 'd2903
      10'd733  : in_data <= 14'h0e93; // 'd3731
      10'd734  : in_data <= 14'h015e; // 'd350
      10'd735  : in_data <= 14'h0de5; // 'd3557
      10'd736  : in_data <= 14'h0072; // 'd114
      10'd737  : in_data <= 14'h0ff9; // 'd4089
      10'd738  : in_data <= 14'h01ab; // 'd427
      10'd739  : in_data <= 14'h00a8; // 'd168
      10'd740  : in_data <= 14'h0b22; // 'd2850
      10'd741  : in_data <= 14'h0f90; // 'd3984
      10'd742  : in_data <= 14'h0796; // 'd1942
      10'd743  : in_data <= 14'h0326; // 'd806
      10'd744  : in_data <= 14'h04c5; // 'd1221
      10'd745  : in_data <= 14'h01f3; // 'd499
      10'd746  : in_data <= 14'h0955; // 'd2389
      10'd747  : in_data <= 14'h0a06; // 'd2566
      10'd748  : in_data <= 14'h0890; // 'd2192
      10'd749  : in_data <= 14'h0325; // 'd805
      10'd750  : in_data <= 14'h00e4; // 'd228
      10'd751  : in_data <= 14'h0373; // 'd883
      10'd752  : in_data <= 14'h02d4; // 'd724
      10'd753  : in_data <= 14'h0b3f; // 'd2879
      10'd754  : in_data <= 14'h0e97; // 'd3735
      10'd755  : in_data <= 14'h016e; // 'd366
      10'd756  : in_data <= 14'h0a5e; // 'd2654
      10'd757  : in_data <= 14'h0456; // 'd1110
      10'd758  : in_data <= 14'h1061; // 'd4193
      10'd759  : in_data <= 14'h054f; // 'd1359
      10'd760  : in_data <= 14'h107b; // 'd4219
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      11'd0    : out_data_ref <= 8'h36;
      11'd1    : out_data_ref <= 8'hc9;
      11'd2    : out_data_ref <= 8'h69;
      11'd3    : out_data_ref <= 8'hcf;
      11'd4    : out_data_ref <= 8'h10;
      11'd5    : out_data_ref <= 8'h08;
      11'd6    : out_data_ref <= 8'ha6;
      11'd7    : out_data_ref <= 8'haa;
      11'd8    : out_data_ref <= 8'h95;
      11'd9    : out_data_ref <= 8'h51;
      11'd10   : out_data_ref <= 8'ha7;
      11'd11   : out_data_ref <= 8'h84;
      11'd12   : out_data_ref <= 8'h94;
      11'd13   : out_data_ref <= 8'h1c;
      11'd14   : out_data_ref <= 8'h65;
      11'd15   : out_data_ref <= 8'ha9;
      11'd16   : out_data_ref <= 8'hbf;
      11'd17   : out_data_ref <= 8'h68;
      11'd18   : out_data_ref <= 8'hc2;
      11'd19   : out_data_ref <= 8'hdc;
      11'd20   : out_data_ref <= 8'h33;
      11'd21   : out_data_ref <= 8'hfa;
      11'd22   : out_data_ref <= 8'h36;
      11'd23   : out_data_ref <= 8'hb5;
      11'd24   : out_data_ref <= 8'hd2;
      11'd25   : out_data_ref <= 8'h66;
      11'd26   : out_data_ref <= 8'hb2;
      11'd27   : out_data_ref <= 8'h51;
      11'd28   : out_data_ref <= 8'h71;
      11'd29   : out_data_ref <= 8'hb3;
      11'd30   : out_data_ref <= 8'h46;
      11'd31   : out_data_ref <= 8'h67;
      11'd32   : out_data_ref <= 8'h9f;
      11'd33   : out_data_ref <= 8'h2d;
      11'd34   : out_data_ref <= 8'h22;
      11'd35   : out_data_ref <= 8'hbf;
      11'd36   : out_data_ref <= 8'h31;
      11'd37   : out_data_ref <= 8'h23;
      11'd38   : out_data_ref <= 8'ha7;
      11'd39   : out_data_ref <= 8'h9c;
      11'd40   : out_data_ref <= 8'h79;
      11'd41   : out_data_ref <= 8'h0d;
      11'd42   : out_data_ref <= 8'h6d;
      11'd43   : out_data_ref <= 8'hec;
      11'd44   : out_data_ref <= 8'h68;
      11'd45   : out_data_ref <= 8'he1;
      11'd46   : out_data_ref <= 8'hbc;
      11'd47   : out_data_ref <= 8'h44;
      11'd48   : out_data_ref <= 8'h42;
      11'd49   : out_data_ref <= 8'h0a;
      11'd50   : out_data_ref <= 8'h68;
      11'd51   : out_data_ref <= 8'h24;
      11'd52   : out_data_ref <= 8'hf5;
      11'd53   : out_data_ref <= 8'h35;
      11'd54   : out_data_ref <= 8'h7c;
      11'd55   : out_data_ref <= 8'h78;
      11'd56   : out_data_ref <= 8'he3;
      11'd57   : out_data_ref <= 8'hc3;
      11'd58   : out_data_ref <= 8'h36;
      11'd59   : out_data_ref <= 8'hfe;
      11'd60   : out_data_ref <= 8'he0;
      11'd61   : out_data_ref <= 8'h55;
      11'd62   : out_data_ref <= 8'h1e;
      11'd63   : out_data_ref <= 8'h62;
      11'd64   : out_data_ref <= 8'h0d;
      11'd65   : out_data_ref <= 8'hcb;
      11'd66   : out_data_ref <= 8'h97;
      11'd67   : out_data_ref <= 8'h5f;
      11'd68   : out_data_ref <= 8'h56;
      11'd69   : out_data_ref <= 8'h36;
      11'd70   : out_data_ref <= 8'h82;
      11'd71   : out_data_ref <= 8'ha3;
      11'd72   : out_data_ref <= 8'h12;
      11'd73   : out_data_ref <= 8'ha3;
      11'd74   : out_data_ref <= 8'h35;
      11'd75   : out_data_ref <= 8'h3b;
      11'd76   : out_data_ref <= 8'h52;
      11'd77   : out_data_ref <= 8'h1c;
      11'd78   : out_data_ref <= 8'h72;
      11'd79   : out_data_ref <= 8'h7f;
      11'd80   : out_data_ref <= 8'h57;
      11'd81   : out_data_ref <= 8'hca;
      11'd82   : out_data_ref <= 8'hbe;
      11'd83   : out_data_ref <= 8'hd0;
      11'd84   : out_data_ref <= 8'hc3;
      11'd85   : out_data_ref <= 8'h22;
      11'd86   : out_data_ref <= 8'h8f;
      11'd87   : out_data_ref <= 8'h09;
      11'd88   : out_data_ref <= 8'h31;
      11'd89   : out_data_ref <= 8'h7c;
      11'd90   : out_data_ref <= 8'hae;
      11'd91   : out_data_ref <= 8'h8b;
      11'd92   : out_data_ref <= 8'h58;
      11'd93   : out_data_ref <= 8'h15;
      11'd94   : out_data_ref <= 8'h8e;
      11'd95   : out_data_ref <= 8'hbf;
      11'd96   : out_data_ref <= 8'h5b;
      11'd97   : out_data_ref <= 8'h26;
      11'd98   : out_data_ref <= 8'hbd;
      11'd99   : out_data_ref <= 8'hc6;
      11'd100  : out_data_ref <= 8'he6;
      11'd101  : out_data_ref <= 8'h36;
      11'd102  : out_data_ref <= 8'h5a;
      11'd103  : out_data_ref <= 8'ha6;
      11'd104  : out_data_ref <= 8'h01;
      11'd105  : out_data_ref <= 8'hac;
      11'd106  : out_data_ref <= 8'had;
      11'd107  : out_data_ref <= 8'h2a;
      11'd108  : out_data_ref <= 8'hbd;
      11'd109  : out_data_ref <= 8'h37;
      11'd110  : out_data_ref <= 8'hf5;
      11'd111  : out_data_ref <= 8'h83;
      11'd112  : out_data_ref <= 8'h0d;
      11'd113  : out_data_ref <= 8'h0b;
      11'd114  : out_data_ref <= 8'hbf;
      11'd115  : out_data_ref <= 8'he3;
      11'd116  : out_data_ref <= 8'h55;
      11'd117  : out_data_ref <= 8'h70;
      11'd118  : out_data_ref <= 8'h5c;
      11'd119  : out_data_ref <= 8'h0a;
      11'd120  : out_data_ref <= 8'h62;
      11'd121  : out_data_ref <= 8'hb7;
      11'd122  : out_data_ref <= 8'h6a;
      11'd123  : out_data_ref <= 8'h5c;
      11'd124  : out_data_ref <= 8'h91;
      11'd125  : out_data_ref <= 8'h0a;
      11'd126  : out_data_ref <= 8'hd0;
      11'd127  : out_data_ref <= 8'h4e;
      11'd128  : out_data_ref <= 8'h55;
      11'd129  : out_data_ref <= 8'he5;
      11'd130  : out_data_ref <= 8'hda;
      11'd131  : out_data_ref <= 8'hd7;
      11'd132  : out_data_ref <= 8'h49;
      11'd133  : out_data_ref <= 8'hc7;
      11'd134  : out_data_ref <= 8'h39;
      11'd135  : out_data_ref <= 8'h3d;
      11'd136  : out_data_ref <= 8'h2e;
      11'd137  : out_data_ref <= 8'h2e;
      11'd138  : out_data_ref <= 8'h8a;
      11'd139  : out_data_ref <= 8'hb6;
      11'd140  : out_data_ref <= 8'h43;
      11'd141  : out_data_ref <= 8'he6;
      11'd142  : out_data_ref <= 8'h2e;
      11'd143  : out_data_ref <= 8'h47;
      11'd144  : out_data_ref <= 8'h57;
      11'd145  : out_data_ref <= 8'had;
      11'd146  : out_data_ref <= 8'h22;
      11'd147  : out_data_ref <= 8'h01;
      11'd148  : out_data_ref <= 8'hca;
      11'd149  : out_data_ref <= 8'ha3;
      11'd150  : out_data_ref <= 8'h32;
      11'd151  : out_data_ref <= 8'h03;
      11'd152  : out_data_ref <= 8'hf5;
      11'd153  : out_data_ref <= 8'h3b;
      11'd154  : out_data_ref <= 8'h4a;
      11'd155  : out_data_ref <= 8'h9d;
      11'd156  : out_data_ref <= 8'h47;
      11'd157  : out_data_ref <= 8'h57;
      11'd158  : out_data_ref <= 8'he7;
      11'd159  : out_data_ref <= 8'h27;
      11'd160  : out_data_ref <= 8'h4d;
      11'd161  : out_data_ref <= 8'h72;
      11'd162  : out_data_ref <= 8'hbd;
      11'd163  : out_data_ref <= 8'hb0;
      11'd164  : out_data_ref <= 8'h36;
      11'd165  : out_data_ref <= 8'ha3;
      11'd166  : out_data_ref <= 8'h1d;
      11'd167  : out_data_ref <= 8'h7d;
      11'd168  : out_data_ref <= 8'he1;
      11'd169  : out_data_ref <= 8'h1e;
      11'd170  : out_data_ref <= 8'h5d;
      11'd171  : out_data_ref <= 8'h1c;
      11'd172  : out_data_ref <= 8'h66;
      11'd173  : out_data_ref <= 8'hcf;
      11'd174  : out_data_ref <= 8'h30;
      11'd175  : out_data_ref <= 8'h59;
      11'd176  : out_data_ref <= 8'hf3;
      11'd177  : out_data_ref <= 8'h3b;
      11'd178  : out_data_ref <= 8'h6a;
      11'd179  : out_data_ref <= 8'h29;
      11'd180  : out_data_ref <= 8'h72;
      11'd181  : out_data_ref <= 8'hc1;
      11'd182  : out_data_ref <= 8'he1;
      11'd183  : out_data_ref <= 8'hd9;
      11'd184  : out_data_ref <= 8'hc9;
      11'd185  : out_data_ref <= 8'hfb;
      11'd186  : out_data_ref <= 8'h2a;
      11'd187  : out_data_ref <= 8'heb;
      11'd188  : out_data_ref <= 8'hc7;
      11'd189  : out_data_ref <= 8'h8b;
      11'd190  : out_data_ref <= 8'h2c;
      11'd191  : out_data_ref <= 8'h05;
      11'd192  : out_data_ref <= 8'h5d;
      11'd193  : out_data_ref <= 8'h48;
      11'd194  : out_data_ref <= 8'hd7;
      11'd195  : out_data_ref <= 8'h9c;
      11'd196  : out_data_ref <= 8'h3a;
      11'd197  : out_data_ref <= 8'h7c;
      11'd198  : out_data_ref <= 8'h99;
      11'd199  : out_data_ref <= 8'h6c;
      11'd200  : out_data_ref <= 8'h08;
      11'd201  : out_data_ref <= 8'hb7;
      11'd202  : out_data_ref <= 8'hde;
      11'd203  : out_data_ref <= 8'hf0;
      11'd204  : out_data_ref <= 8'h79;
      11'd205  : out_data_ref <= 8'h1c;
      11'd206  : out_data_ref <= 8'hde;
      11'd207  : out_data_ref <= 8'h89;
      11'd208  : out_data_ref <= 8'h50;
      11'd209  : out_data_ref <= 8'h53;
      11'd210  : out_data_ref <= 8'h88;
      11'd211  : out_data_ref <= 8'h5d;
      11'd212  : out_data_ref <= 8'h8d;
      11'd213  : out_data_ref <= 8'ha1;
      11'd214  : out_data_ref <= 8'hd2;
      11'd215  : out_data_ref <= 8'h54;
      11'd216  : out_data_ref <= 8'hee;
      11'd217  : out_data_ref <= 8'h19;
      11'd218  : out_data_ref <= 8'hc0;
      11'd219  : out_data_ref <= 8'h90;
      11'd220  : out_data_ref <= 8'haf;
      11'd221  : out_data_ref <= 8'h34;
      11'd222  : out_data_ref <= 8'hf4;
      11'd223  : out_data_ref <= 8'h72;
      11'd224  : out_data_ref <= 8'h0b;
      11'd225  : out_data_ref <= 8'h0b;
      11'd226  : out_data_ref <= 8'h77;
      11'd227  : out_data_ref <= 8'h13;
      11'd228  : out_data_ref <= 8'h91;
      11'd229  : out_data_ref <= 8'h08;
      11'd230  : out_data_ref <= 8'hd8;
      11'd231  : out_data_ref <= 8'h49;
      11'd232  : out_data_ref <= 8'h89;
      11'd233  : out_data_ref <= 8'h82;
      11'd234  : out_data_ref <= 8'hfe;
      11'd235  : out_data_ref <= 8'hab;
      11'd236  : out_data_ref <= 8'h0b;
      11'd237  : out_data_ref <= 8'h54;
      11'd238  : out_data_ref <= 8'h93;
      11'd239  : out_data_ref <= 8'h4c;
      11'd240  : out_data_ref <= 8'hee;
      11'd241  : out_data_ref <= 8'h3d;
      11'd242  : out_data_ref <= 8'hcd;
      11'd243  : out_data_ref <= 8'h24;
      11'd244  : out_data_ref <= 8'hb0;
      11'd245  : out_data_ref <= 8'h49;
      11'd246  : out_data_ref <= 8'hf9;
      11'd247  : out_data_ref <= 8'h81;
      11'd248  : out_data_ref <= 8'ha8;
      11'd249  : out_data_ref <= 8'h4c;
      11'd250  : out_data_ref <= 8'h92;
      11'd251  : out_data_ref <= 8'h80;
      11'd252  : out_data_ref <= 8'h28;
      11'd253  : out_data_ref <= 8'ha6;
      11'd254  : out_data_ref <= 8'h4a;
      11'd255  : out_data_ref <= 8'h26;
      11'd256  : out_data_ref <= 8'hcd;
      11'd257  : out_data_ref <= 8'hf8;
      11'd258  : out_data_ref <= 8'h70;
      11'd259  : out_data_ref <= 8'h52;
      11'd260  : out_data_ref <= 8'h31;
      11'd261  : out_data_ref <= 8'h3c;
      11'd262  : out_data_ref <= 8'h3e;
      11'd263  : out_data_ref <= 8'h50;
      11'd264  : out_data_ref <= 8'hb2;
      11'd265  : out_data_ref <= 8'he1;
      11'd266  : out_data_ref <= 8'hf5;
      11'd267  : out_data_ref <= 8'h39;
      11'd268  : out_data_ref <= 8'h39;
      11'd269  : out_data_ref <= 8'h45;
      11'd270  : out_data_ref <= 8'h02;
      11'd271  : out_data_ref <= 8'h43;
      11'd272  : out_data_ref <= 8'h3c;
      11'd273  : out_data_ref <= 8'h09;
      11'd274  : out_data_ref <= 8'h62;
      11'd275  : out_data_ref <= 8'h99;
      11'd276  : out_data_ref <= 8'h6c;
      11'd277  : out_data_ref <= 8'h35;
      11'd278  : out_data_ref <= 8'h99;
      11'd279  : out_data_ref <= 8'h18;
      11'd280  : out_data_ref <= 8'h9b;
      11'd281  : out_data_ref <= 8'h15;
      11'd282  : out_data_ref <= 8'h17;
      11'd283  : out_data_ref <= 8'h42;
      11'd284  : out_data_ref <= 8'h81;
      11'd285  : out_data_ref <= 8'hb6;
      11'd286  : out_data_ref <= 8'h59;
      11'd287  : out_data_ref <= 8'h5b;
      11'd288  : out_data_ref <= 8'h56;
      11'd289  : out_data_ref <= 8'h7b;
      11'd290  : out_data_ref <= 8'h8c;
      11'd291  : out_data_ref <= 8'h4c;
      11'd292  : out_data_ref <= 8'hd8;
      11'd293  : out_data_ref <= 8'h09;
      11'd294  : out_data_ref <= 8'h02;
      11'd295  : out_data_ref <= 8'h86;
      11'd296  : out_data_ref <= 8'h0e;
      11'd297  : out_data_ref <= 8'h61;
      11'd298  : out_data_ref <= 8'h3a;
      11'd299  : out_data_ref <= 8'he1;
      11'd300  : out_data_ref <= 8'h90;
      11'd301  : out_data_ref <= 8'h6a;
      11'd302  : out_data_ref <= 8'h55;
      11'd303  : out_data_ref <= 8'h60;
      11'd304  : out_data_ref <= 8'h7c;
      11'd305  : out_data_ref <= 8'hbf;
      11'd306  : out_data_ref <= 8'h0e;
      11'd307  : out_data_ref <= 8'h11;
      11'd308  : out_data_ref <= 8'had;
      11'd309  : out_data_ref <= 8'h6c;
      11'd310  : out_data_ref <= 8'h0c;
      11'd311  : out_data_ref <= 8'h0d;
      11'd312  : out_data_ref <= 8'hf3;
      11'd313  : out_data_ref <= 8'h8c;
      11'd314  : out_data_ref <= 8'h00;
      11'd315  : out_data_ref <= 8'h6a;
      11'd316  : out_data_ref <= 8'h5f;
      11'd317  : out_data_ref <= 8'h53;
      11'd318  : out_data_ref <= 8'h5f;
      11'd319  : out_data_ref <= 8'ha6;
      11'd320  : out_data_ref <= 8'he6;
      11'd321  : out_data_ref <= 8'hfb;
      11'd322  : out_data_ref <= 8'h49;
      11'd323  : out_data_ref <= 8'hd1;
      11'd324  : out_data_ref <= 8'h0b;
      11'd325  : out_data_ref <= 8'h78;
      11'd326  : out_data_ref <= 8'hb9;
      11'd327  : out_data_ref <= 8'hcb;
      11'd328  : out_data_ref <= 8'h64;
      11'd329  : out_data_ref <= 8'h73;
      11'd330  : out_data_ref <= 8'hbf;
      11'd331  : out_data_ref <= 8'h06;
      11'd332  : out_data_ref <= 8'h30;
      11'd333  : out_data_ref <= 8'h51;
      11'd334  : out_data_ref <= 8'h8d;
      11'd335  : out_data_ref <= 8'hb6;
      11'd336  : out_data_ref <= 8'hfd;
      11'd337  : out_data_ref <= 8'hec;
      11'd338  : out_data_ref <= 8'hfd;
      11'd339  : out_data_ref <= 8'h70;
      11'd340  : out_data_ref <= 8'hde;
      11'd341  : out_data_ref <= 8'hd2;
      11'd342  : out_data_ref <= 8'h01;
      11'd343  : out_data_ref <= 8'hc7;
      11'd344  : out_data_ref <= 8'he3;
      11'd345  : out_data_ref <= 8'h5f;
      11'd346  : out_data_ref <= 8'hfb;
      11'd347  : out_data_ref <= 8'h3b;
      11'd348  : out_data_ref <= 8'hb7;
      11'd349  : out_data_ref <= 8'h8d;
      11'd350  : out_data_ref <= 8'h8a;
      11'd351  : out_data_ref <= 8'hec;
      11'd352  : out_data_ref <= 8'h18;
      11'd353  : out_data_ref <= 8'h1f;
      11'd354  : out_data_ref <= 8'h6d;
      11'd355  : out_data_ref <= 8'he9;
      11'd356  : out_data_ref <= 8'h60;
      11'd357  : out_data_ref <= 8'hc3;
      11'd358  : out_data_ref <= 8'h16;
      11'd359  : out_data_ref <= 8'hfe;
      11'd360  : out_data_ref <= 8'h35;
      11'd361  : out_data_ref <= 8'h4b;
      11'd362  : out_data_ref <= 8'h7c;
      11'd363  : out_data_ref <= 8'hc6;
      11'd364  : out_data_ref <= 8'h9e;
      11'd365  : out_data_ref <= 8'h80;
      11'd366  : out_data_ref <= 8'h48;
      11'd367  : out_data_ref <= 8'h20;
      11'd368  : out_data_ref <= 8'h19;
      11'd369  : out_data_ref <= 8'h65;
      11'd370  : out_data_ref <= 8'haa;
      11'd371  : out_data_ref <= 8'hfe;
      11'd372  : out_data_ref <= 8'hf4;
      11'd373  : out_data_ref <= 8'hea;
      11'd374  : out_data_ref <= 8'h3f;
      11'd375  : out_data_ref <= 8'h80;
      11'd376  : out_data_ref <= 8'h87;
      11'd377  : out_data_ref <= 8'h37;
      11'd378  : out_data_ref <= 8'hff;
      11'd379  : out_data_ref <= 8'h45;
      11'd380  : out_data_ref <= 8'h25;
      11'd381  : out_data_ref <= 8'h5a;
      11'd382  : out_data_ref <= 8'h17;
      11'd383  : out_data_ref <= 8'h79;
      11'd384  : out_data_ref <= 8'hde;
      11'd385  : out_data_ref <= 8'h57;
      11'd386  : out_data_ref <= 8'ha4;
      11'd387  : out_data_ref <= 8'hb6;
      11'd388  : out_data_ref <= 8'h8d;
      11'd389  : out_data_ref <= 8'hb5;
      11'd390  : out_data_ref <= 8'h87;
      11'd391  : out_data_ref <= 8'h26;
      11'd392  : out_data_ref <= 8'h3d;
      11'd393  : out_data_ref <= 8'h7b;
      11'd394  : out_data_ref <= 8'h7f;
      11'd395  : out_data_ref <= 8'h6c;
      11'd396  : out_data_ref <= 8'hb0;
      11'd397  : out_data_ref <= 8'h7d;
      11'd398  : out_data_ref <= 8'h8b;
      11'd399  : out_data_ref <= 8'h01;
      11'd400  : out_data_ref <= 8'h22;
      11'd401  : out_data_ref <= 8'h4d;
      11'd402  : out_data_ref <= 8'hd2;
      11'd403  : out_data_ref <= 8'h91;
      11'd404  : out_data_ref <= 8'h23;
      11'd405  : out_data_ref <= 8'h7e;
      11'd406  : out_data_ref <= 8'hfd;
      11'd407  : out_data_ref <= 8'h9c;
      11'd408  : out_data_ref <= 8'h01;
      11'd409  : out_data_ref <= 8'h67;
      11'd410  : out_data_ref <= 8'h6e;
      11'd411  : out_data_ref <= 8'h30;
      11'd412  : out_data_ref <= 8'h15;
      11'd413  : out_data_ref <= 8'h4a;
      11'd414  : out_data_ref <= 8'h2a;
      11'd415  : out_data_ref <= 8'h7d;
      11'd416  : out_data_ref <= 8'h60;
      11'd417  : out_data_ref <= 8'h17;
      11'd418  : out_data_ref <= 8'h45;
      11'd419  : out_data_ref <= 8'h36;
      11'd420  : out_data_ref <= 8'h58;
      11'd421  : out_data_ref <= 8'h0f;
      11'd422  : out_data_ref <= 8'he6;
      11'd423  : out_data_ref <= 8'h4e;
      11'd424  : out_data_ref <= 8'hfe;
      11'd425  : out_data_ref <= 8'hdd;
      11'd426  : out_data_ref <= 8'ha5;
      11'd427  : out_data_ref <= 8'hfb;
      11'd428  : out_data_ref <= 8'h42;
      11'd429  : out_data_ref <= 8'hc1;
      11'd430  : out_data_ref <= 8'h3e;
      11'd431  : out_data_ref <= 8'hd8;
      11'd432  : out_data_ref <= 8'hc5;
      11'd433  : out_data_ref <= 8'h76;
      11'd434  : out_data_ref <= 8'h8a;
      11'd435  : out_data_ref <= 8'h3c;
      11'd436  : out_data_ref <= 8'hbc;
      11'd437  : out_data_ref <= 8'hae;
      11'd438  : out_data_ref <= 8'h7a;
      11'd439  : out_data_ref <= 8'h23;
      11'd440  : out_data_ref <= 8'h43;
      11'd441  : out_data_ref <= 8'hb3;
      11'd442  : out_data_ref <= 8'h12;
      11'd443  : out_data_ref <= 8'h8c;
      11'd444  : out_data_ref <= 8'hd5;
      11'd445  : out_data_ref <= 8'hc1;
      11'd446  : out_data_ref <= 8'hc6;
      11'd447  : out_data_ref <= 8'h63;
      11'd448  : out_data_ref <= 8'ha0;
      11'd449  : out_data_ref <= 8'h7c;
      11'd450  : out_data_ref <= 8'h7d;
      11'd451  : out_data_ref <= 8'hc0;
      11'd452  : out_data_ref <= 8'he1;
      11'd453  : out_data_ref <= 8'he2;
      11'd454  : out_data_ref <= 8'h64;
      11'd455  : out_data_ref <= 8'h2c;
      11'd456  : out_data_ref <= 8'h0d;
      11'd457  : out_data_ref <= 8'h9a;
      11'd458  : out_data_ref <= 8'h02;
      11'd459  : out_data_ref <= 8'hf3;
      11'd460  : out_data_ref <= 8'h49;
      11'd461  : out_data_ref <= 8'hc9;
      11'd462  : out_data_ref <= 8'h64;
      11'd463  : out_data_ref <= 8'h15;
      11'd464  : out_data_ref <= 8'h4a;
      11'd465  : out_data_ref <= 8'h6c;
      11'd466  : out_data_ref <= 8'h43;
      11'd467  : out_data_ref <= 8'h08;
      11'd468  : out_data_ref <= 8'hd8;
      11'd469  : out_data_ref <= 8'hec;
      11'd470  : out_data_ref <= 8'hf3;
      11'd471  : out_data_ref <= 8'h0f;
      11'd472  : out_data_ref <= 8'h47;
      11'd473  : out_data_ref <= 8'he9;
      11'd474  : out_data_ref <= 8'ha8;
      11'd475  : out_data_ref <= 8'h1e;
      11'd476  : out_data_ref <= 8'hed;
      11'd477  : out_data_ref <= 8'h2a;
      11'd478  : out_data_ref <= 8'h32;
      11'd479  : out_data_ref <= 8'ha2;
      11'd480  : out_data_ref <= 8'hbb;
      11'd481  : out_data_ref <= 8'h44;
      11'd482  : out_data_ref <= 8'hdf;
      11'd483  : out_data_ref <= 8'hc3;
      11'd484  : out_data_ref <= 8'h6a;
      11'd485  : out_data_ref <= 8'h28;
      11'd486  : out_data_ref <= 8'ha6;
      11'd487  : out_data_ref <= 8'h6a;
      11'd488  : out_data_ref <= 8'he7;
      11'd489  : out_data_ref <= 8'h7b;
      11'd490  : out_data_ref <= 8'hb1;
      11'd491  : out_data_ref <= 8'h39;
      11'd492  : out_data_ref <= 8'hfa;
      11'd493  : out_data_ref <= 8'h41;
      11'd494  : out_data_ref <= 8'h6b;
      11'd495  : out_data_ref <= 8'h63;
      11'd496  : out_data_ref <= 8'h27;
      11'd497  : out_data_ref <= 8'hee;
      11'd498  : out_data_ref <= 8'hfe;
      11'd499  : out_data_ref <= 8'h33;
      11'd500  : out_data_ref <= 8'h63;
      11'd501  : out_data_ref <= 8'h24;
      11'd502  : out_data_ref <= 8'h69;
      11'd503  : out_data_ref <= 8'hcc;
      11'd504  : out_data_ref <= 8'hc2;
      11'd505  : out_data_ref <= 8'h12;
      11'd506  : out_data_ref <= 8'h29;
      11'd507  : out_data_ref <= 8'h58;
      11'd508  : out_data_ref <= 8'h75;
      11'd509  : out_data_ref <= 8'h73;
      11'd510  : out_data_ref <= 8'hc4;
      11'd511  : out_data_ref <= 8'hf7;
      11'd512  : out_data_ref <= 8'h75;
      11'd513  : out_data_ref <= 8'h2c;
      11'd514  : out_data_ref <= 8'he1;
      11'd515  : out_data_ref <= 8'hcc;
      11'd516  : out_data_ref <= 8'h79;
      11'd517  : out_data_ref <= 8'hca;
      11'd518  : out_data_ref <= 8'h0c;
      11'd519  : out_data_ref <= 8'h6b;
      11'd520  : out_data_ref <= 8'hda;
      11'd521  : out_data_ref <= 8'h08;
      11'd522  : out_data_ref <= 8'hcd;
      11'd523  : out_data_ref <= 8'h79;
      11'd524  : out_data_ref <= 8'he2;
      11'd525  : out_data_ref <= 8'h57;
      11'd526  : out_data_ref <= 8'h20;
      11'd527  : out_data_ref <= 8'hd2;
      11'd528  : out_data_ref <= 8'hd9;
      11'd529  : out_data_ref <= 8'h09;
      11'd530  : out_data_ref <= 8'h2e;
      11'd531  : out_data_ref <= 8'ha2;
      11'd532  : out_data_ref <= 8'hab;
      11'd533  : out_data_ref <= 8'h13;
      11'd534  : out_data_ref <= 8'hf3;
      11'd535  : out_data_ref <= 8'h1e;
      11'd536  : out_data_ref <= 8'h9a;
      11'd537  : out_data_ref <= 8'h3a;
      11'd538  : out_data_ref <= 8'hf1;
      11'd539  : out_data_ref <= 8'hc6;
      11'd540  : out_data_ref <= 8'h9f;
      11'd541  : out_data_ref <= 8'hc6;
      11'd542  : out_data_ref <= 8'h37;
      11'd543  : out_data_ref <= 8'h9d;
      11'd544  : out_data_ref <= 8'h8e;
      11'd545  : out_data_ref <= 8'h2a;
      11'd546  : out_data_ref <= 8'hd2;
      11'd547  : out_data_ref <= 8'hb8;
      11'd548  : out_data_ref <= 8'h7b;
      11'd549  : out_data_ref <= 8'h51;
      11'd550  : out_data_ref <= 8'h4c;
      11'd551  : out_data_ref <= 8'h81;
      11'd552  : out_data_ref <= 8'h7a;
      11'd553  : out_data_ref <= 8'h08;
      11'd554  : out_data_ref <= 8'h73;
      11'd555  : out_data_ref <= 8'h38;
      11'd556  : out_data_ref <= 8'hb7;
      11'd557  : out_data_ref <= 8'hb0;
      11'd558  : out_data_ref <= 8'h73;
      11'd559  : out_data_ref <= 8'h6b;
      11'd560  : out_data_ref <= 8'h89;
      11'd561  : out_data_ref <= 8'h54;
      11'd562  : out_data_ref <= 8'hde;
      11'd563  : out_data_ref <= 8'h92;
      11'd564  : out_data_ref <= 8'h23;
      11'd565  : out_data_ref <= 8'h22;
      11'd566  : out_data_ref <= 8'h5b;
      11'd567  : out_data_ref <= 8'h40;
      11'd568  : out_data_ref <= 8'h07;
      11'd569  : out_data_ref <= 8'h9c;
      11'd570  : out_data_ref <= 8'h92;
      11'd571  : out_data_ref <= 8'h60;
      11'd572  : out_data_ref <= 8'h12;
      11'd573  : out_data_ref <= 8'h48;
      11'd574  : out_data_ref <= 8'hc1;
      11'd575  : out_data_ref <= 8'h4b;
      11'd576  : out_data_ref <= 8'h21;
      11'd577  : out_data_ref <= 8'h04;
      11'd578  : out_data_ref <= 8'h90;
      11'd579  : out_data_ref <= 8'h1e;
      11'd580  : out_data_ref <= 8'h74;
      11'd581  : out_data_ref <= 8'hf8;
      11'd582  : out_data_ref <= 8'h49;
      11'd583  : out_data_ref <= 8'hd9;
      11'd584  : out_data_ref <= 8'hee;
      11'd585  : out_data_ref <= 8'he9;
      11'd586  : out_data_ref <= 8'hf5;
      11'd587  : out_data_ref <= 8'h63;
      11'd588  : out_data_ref <= 8'h6c;
      11'd589  : out_data_ref <= 8'h1d;
      11'd590  : out_data_ref <= 8'had;
      11'd591  : out_data_ref <= 8'h60;
      11'd592  : out_data_ref <= 8'h31;
      11'd593  : out_data_ref <= 8'hab;
      11'd594  : out_data_ref <= 8'h47;
      11'd595  : out_data_ref <= 8'h7c;
      11'd596  : out_data_ref <= 8'h57;
      11'd597  : out_data_ref <= 8'h31;
      11'd598  : out_data_ref <= 8'h97;
      11'd599  : out_data_ref <= 8'he7;
      11'd600  : out_data_ref <= 8'heb;
      11'd601  : out_data_ref <= 8'h6c;
      11'd602  : out_data_ref <= 8'he5;
      11'd603  : out_data_ref <= 8'h35;
      11'd604  : out_data_ref <= 8'hd9;
      11'd605  : out_data_ref <= 8'hf0;
      11'd606  : out_data_ref <= 8'hf6;
      11'd607  : out_data_ref <= 8'h91;
      11'd608  : out_data_ref <= 8'h83;
      11'd609  : out_data_ref <= 8'hdd;
      11'd610  : out_data_ref <= 8'h9d;
      11'd611  : out_data_ref <= 8'hf5;
      11'd612  : out_data_ref <= 8'h52;
      11'd613  : out_data_ref <= 8'h15;
      11'd614  : out_data_ref <= 8'h95;
      11'd615  : out_data_ref <= 8'he5;
      11'd616  : out_data_ref <= 8'hc9;
      11'd617  : out_data_ref <= 8'he9;
      11'd618  : out_data_ref <= 8'h8d;
      11'd619  : out_data_ref <= 8'h84;
      11'd620  : out_data_ref <= 8'h6c;
      11'd621  : out_data_ref <= 8'he0;
      11'd622  : out_data_ref <= 8'h8a;
      11'd623  : out_data_ref <= 8'ha6;
      11'd624  : out_data_ref <= 8'h55;
      11'd625  : out_data_ref <= 8'hb7;
      11'd626  : out_data_ref <= 8'h0c;
      11'd627  : out_data_ref <= 8'hc0;
      11'd628  : out_data_ref <= 8'hd8;
      11'd629  : out_data_ref <= 8'h04;
      11'd630  : out_data_ref <= 8'h14;
      11'd631  : out_data_ref <= 8'h01;
      11'd632  : out_data_ref <= 8'h92;
      11'd633  : out_data_ref <= 8'h96;
      11'd634  : out_data_ref <= 8'h90;
      11'd635  : out_data_ref <= 8'h29;
      11'd636  : out_data_ref <= 8'h8f;
      11'd637  : out_data_ref <= 8'h64;
      11'd638  : out_data_ref <= 8'h5d;
      11'd639  : out_data_ref <= 8'h91;
      11'd640  : out_data_ref <= 8'h12;
      11'd641  : out_data_ref <= 8'hdb;
      11'd642  : out_data_ref <= 8'hb0;
      11'd643  : out_data_ref <= 8'h3b;
      11'd644  : out_data_ref <= 8'h18;
      11'd645  : out_data_ref <= 8'h9c;
      11'd646  : out_data_ref <= 8'hdb;
      11'd647  : out_data_ref <= 8'h1f;
      11'd648  : out_data_ref <= 8'hcf;
      11'd649  : out_data_ref <= 8'h4d;
      11'd650  : out_data_ref <= 8'h51;
      11'd651  : out_data_ref <= 8'h2f;
      11'd652  : out_data_ref <= 8'h68;
      11'd653  : out_data_ref <= 8'h74;
      11'd654  : out_data_ref <= 8'hb4;
      11'd655  : out_data_ref <= 8'h09;
      11'd656  : out_data_ref <= 8'hbf;
      11'd657  : out_data_ref <= 8'h55;
      11'd658  : out_data_ref <= 8'hee;
      11'd659  : out_data_ref <= 8'h1c;
      11'd660  : out_data_ref <= 8'hc2;
      11'd661  : out_data_ref <= 8'h84;
      11'd662  : out_data_ref <= 8'ha0;
      11'd663  : out_data_ref <= 8'h5b;
      11'd664  : out_data_ref <= 8'h69;
      11'd665  : out_data_ref <= 8'h8b;
      11'd666  : out_data_ref <= 8'h88;
      11'd667  : out_data_ref <= 8'h18;
      11'd668  : out_data_ref <= 8'hf0;
      11'd669  : out_data_ref <= 8'h43;
      11'd670  : out_data_ref <= 8'hc2;
      11'd671  : out_data_ref <= 8'h59;
      11'd672  : out_data_ref <= 8'h1c;
      11'd673  : out_data_ref <= 8'h9f;
      11'd674  : out_data_ref <= 8'h4a;
      11'd675  : out_data_ref <= 8'hba;
      11'd676  : out_data_ref <= 8'h29;
      11'd677  : out_data_ref <= 8'hcf;
      11'd678  : out_data_ref <= 8'h42;
      11'd679  : out_data_ref <= 8'h59;
      11'd680  : out_data_ref <= 8'h91;
      11'd681  : out_data_ref <= 8'h5d;
      11'd682  : out_data_ref <= 8'h6a;
      11'd683  : out_data_ref <= 8'h0b;
      11'd684  : out_data_ref <= 8'he7;
      11'd685  : out_data_ref <= 8'h1b;
      11'd686  : out_data_ref <= 8'h6b;
      11'd687  : out_data_ref <= 8'h93;
      11'd688  : out_data_ref <= 8'h96;
      11'd689  : out_data_ref <= 8'h3c;
      11'd690  : out_data_ref <= 8'h61;
      11'd691  : out_data_ref <= 8'h8c;
      11'd692  : out_data_ref <= 8'hbb;
      11'd693  : out_data_ref <= 8'h56;
      11'd694  : out_data_ref <= 8'h78;
      11'd695  : out_data_ref <= 8'h38;
      11'd696  : out_data_ref <= 8'he5;
      11'd697  : out_data_ref <= 8'hea;
      11'd698  : out_data_ref <= 8'hde;
      11'd699  : out_data_ref <= 8'h65;
      11'd700  : out_data_ref <= 8'h00;
      11'd701  : out_data_ref <= 8'hde;
      11'd702  : out_data_ref <= 8'h9a;
      11'd703  : out_data_ref <= 8'hd2;
      11'd704  : out_data_ref <= 8'h50;
      11'd705  : out_data_ref <= 8'h08;
      11'd706  : out_data_ref <= 8'h3a;
      11'd707  : out_data_ref <= 8'h01;
      11'd708  : out_data_ref <= 8'heb;
      11'd709  : out_data_ref <= 8'h3e;
      11'd710  : out_data_ref <= 8'hb4;
      11'd711  : out_data_ref <= 8'h4c;
      11'd712  : out_data_ref <= 8'h00;
      11'd713  : out_data_ref <= 8'hee;
      11'd714  : out_data_ref <= 8'hcb;
      11'd715  : out_data_ref <= 8'h2b;
      11'd716  : out_data_ref <= 8'h0f;
      11'd717  : out_data_ref <= 8'h87;
      11'd718  : out_data_ref <= 8'h4c;
      11'd719  : out_data_ref <= 8'hda;
      11'd720  : out_data_ref <= 8'h16;
      11'd721  : out_data_ref <= 8'h5f;
      11'd722  : out_data_ref <= 8'haa;
      11'd723  : out_data_ref <= 8'h65;
      11'd724  : out_data_ref <= 8'h24;
      11'd725  : out_data_ref <= 8'hca;
      11'd726  : out_data_ref <= 8'h13;
      11'd727  : out_data_ref <= 8'hd4;
      11'd728  : out_data_ref <= 8'h35;
      11'd729  : out_data_ref <= 8'hc9;
      11'd730  : out_data_ref <= 8'h38;
      11'd731  : out_data_ref <= 8'hdb;
      11'd732  : out_data_ref <= 8'h94;
      11'd733  : out_data_ref <= 8'h69;
      11'd734  : out_data_ref <= 8'h29;
      11'd735  : out_data_ref <= 8'h2f;
      11'd736  : out_data_ref <= 8'he9;
      11'd737  : out_data_ref <= 8'h72;
      11'd738  : out_data_ref <= 8'h83;
      11'd739  : out_data_ref <= 8'hc6;
      11'd740  : out_data_ref <= 8'h92;
      11'd741  : out_data_ref <= 8'h22;
      11'd742  : out_data_ref <= 8'h10;
      11'd743  : out_data_ref <= 8'h7e;
      11'd744  : out_data_ref <= 8'ha2;
      11'd745  : out_data_ref <= 8'hf9;
      11'd746  : out_data_ref <= 8'hef;
      11'd747  : out_data_ref <= 8'hca;
      11'd748  : out_data_ref <= 8'h1b;
      11'd749  : out_data_ref <= 8'h6d;
      11'd750  : out_data_ref <= 8'h41;
      11'd751  : out_data_ref <= 8'hdc;
      11'd752  : out_data_ref <= 8'ha5;
      11'd753  : out_data_ref <= 8'hb1;
      11'd754  : out_data_ref <= 8'h49;
      11'd755  : out_data_ref <= 8'hb2;
      11'd756  : out_data_ref <= 8'ha8;
      11'd757  : out_data_ref <= 8'hcc;
      11'd758  : out_data_ref <= 8'h22;
      11'd759  : out_data_ref <= 8'h44;
      11'd760  : out_data_ref <= 8'ha1;
      11'd761  : out_data_ref <= 8'hbc;
      11'd762  : out_data_ref <= 8'h54;
      11'd763  : out_data_ref <= 8'h26;
      11'd764  : out_data_ref <= 8'h1c;
      11'd765  : out_data_ref <= 8'hc1;
      11'd766  : out_data_ref <= 8'h17;
      11'd767  : out_data_ref <= 8'h42;
      11'd768  : out_data_ref <= 8'hac;
      11'd769  : out_data_ref <= 8'hd2;
      11'd770  : out_data_ref <= 8'h7b;
      11'd771  : out_data_ref <= 8'h7f;
      11'd772  : out_data_ref <= 8'h23;
      11'd773  : out_data_ref <= 8'h52;
      11'd774  : out_data_ref <= 8'hc3;
      11'd775  : out_data_ref <= 8'h3f;
      11'd776  : out_data_ref <= 8'hb8;
      11'd777  : out_data_ref <= 8'h3f;
      11'd778  : out_data_ref <= 8'he1;
      11'd779  : out_data_ref <= 8'h43;
      11'd780  : out_data_ref <= 8'h38;
      11'd781  : out_data_ref <= 8'h64;
      11'd782  : out_data_ref <= 8'h79;
      11'd783  : out_data_ref <= 8'hd7;
      11'd784  : out_data_ref <= 8'h8d;
      11'd785  : out_data_ref <= 8'h6d;
      11'd786  : out_data_ref <= 8'h5c;
      11'd787  : out_data_ref <= 8'h3e;
      11'd788  : out_data_ref <= 8'h51;
      11'd789  : out_data_ref <= 8'h68;
      11'd790  : out_data_ref <= 8'h4b;
      11'd791  : out_data_ref <= 8'h60;
      11'd792  : out_data_ref <= 8'ha5;
      11'd793  : out_data_ref <= 8'h67;
      11'd794  : out_data_ref <= 8'h14;
      11'd795  : out_data_ref <= 8'h18;
      11'd796  : out_data_ref <= 8'h24;
      11'd797  : out_data_ref <= 8'h49;
      11'd798  : out_data_ref <= 8'hc9;
      11'd799  : out_data_ref <= 8'h43;
      11'd800  : out_data_ref <= 8'h27;
      11'd801  : out_data_ref <= 8'h13;
      11'd802  : out_data_ref <= 8'h9b;
      11'd803  : out_data_ref <= 8'h02;
      11'd804  : out_data_ref <= 8'h89;
      11'd805  : out_data_ref <= 8'hb9;
      11'd806  : out_data_ref <= 8'hbd;
      11'd807  : out_data_ref <= 8'he0;
      11'd808  : out_data_ref <= 8'hae;
      11'd809  : out_data_ref <= 8'h3f;
      11'd810  : out_data_ref <= 8'hef;
      11'd811  : out_data_ref <= 8'h31;
      11'd812  : out_data_ref <= 8'h9f;
      11'd813  : out_data_ref <= 8'he2;
      11'd814  : out_data_ref <= 8'hc6;
      11'd815  : out_data_ref <= 8'h05;
      11'd816  : out_data_ref <= 8'hab;
      11'd817  : out_data_ref <= 8'h55;
      11'd818  : out_data_ref <= 8'h07;
      11'd819  : out_data_ref <= 8'hc8;
      11'd820  : out_data_ref <= 8'h94;
      11'd821  : out_data_ref <= 8'hd2;
      11'd822  : out_data_ref <= 8'hc2;
      11'd823  : out_data_ref <= 8'h76;
      11'd824  : out_data_ref <= 8'h1a;
      11'd825  : out_data_ref <= 8'h3b;
      11'd826  : out_data_ref <= 8'hd3;
      11'd827  : out_data_ref <= 8'hea;
      11'd828  : out_data_ref <= 8'h30;
      11'd829  : out_data_ref <= 8'hf4;
      11'd830  : out_data_ref <= 8'hba;
      11'd831  : out_data_ref <= 8'h92;
      11'd832  : out_data_ref <= 8'h8f;
      11'd833  : out_data_ref <= 8'h9f;
      11'd834  : out_data_ref <= 8'h23;
      11'd835  : out_data_ref <= 8'h30;
      11'd836  : out_data_ref <= 8'h30;
      11'd837  : out_data_ref <= 8'h61;
      11'd838  : out_data_ref <= 8'h61;
      11'd839  : out_data_ref <= 8'h7e;
      11'd840  : out_data_ref <= 8'h2f;
      11'd841  : out_data_ref <= 8'h04;
      11'd842  : out_data_ref <= 8'h2d;
      11'd843  : out_data_ref <= 8'hcf;
      11'd844  : out_data_ref <= 8'h22;
      11'd845  : out_data_ref <= 8'h9a;
      11'd846  : out_data_ref <= 8'hff;
      11'd847  : out_data_ref <= 8'h2c;
      11'd848  : out_data_ref <= 8'h93;
      11'd849  : out_data_ref <= 8'h45;
      11'd850  : out_data_ref <= 8'ha6;
      11'd851  : out_data_ref <= 8'hb3;
      11'd852  : out_data_ref <= 8'hcd;
      11'd853  : out_data_ref <= 8'hcf;
      11'd854  : out_data_ref <= 8'h90;
      11'd855  : out_data_ref <= 8'hd3;
      11'd856  : out_data_ref <= 8'he3;
      11'd857  : out_data_ref <= 8'hbc;
      11'd858  : out_data_ref <= 8'hc3;
      11'd859  : out_data_ref <= 8'ha1;
      11'd860  : out_data_ref <= 8'h11;
      11'd861  : out_data_ref <= 8'h0c;
      11'd862  : out_data_ref <= 8'h85;
      11'd863  : out_data_ref <= 8'h61;
      11'd864  : out_data_ref <= 8'h6b;
      11'd865  : out_data_ref <= 8'hd5;
      11'd866  : out_data_ref <= 8'h85;
      11'd867  : out_data_ref <= 8'hc3;
      11'd868  : out_data_ref <= 8'h1c;
      11'd869  : out_data_ref <= 8'hde;
      11'd870  : out_data_ref <= 8'h3e;
      11'd871  : out_data_ref <= 8'h69;
      11'd872  : out_data_ref <= 8'had;
      11'd873  : out_data_ref <= 8'hc1;
      11'd874  : out_data_ref <= 8'h2a;
      11'd875  : out_data_ref <= 8'h18;
      11'd876  : out_data_ref <= 8'hbf;
      11'd877  : out_data_ref <= 8'ha5;
      11'd878  : out_data_ref <= 8'h79;
      11'd879  : out_data_ref <= 8'h7d;
      11'd880  : out_data_ref <= 8'hf0;
      11'd881  : out_data_ref <= 8'h54;
      11'd882  : out_data_ref <= 8'h34;
      11'd883  : out_data_ref <= 8'h35;
      11'd884  : out_data_ref <= 8'ha7;
      11'd885  : out_data_ref <= 8'hc8;
      11'd886  : out_data_ref <= 8'h74;
      11'd887  : out_data_ref <= 8'ha8;
      11'd888  : out_data_ref <= 8'hac;
      11'd889  : out_data_ref <= 8'hf3;
      11'd890  : out_data_ref <= 8'h78;
      11'd891  : out_data_ref <= 8'h6f;
      11'd892  : out_data_ref <= 8'hcc;
      11'd893  : out_data_ref <= 8'hba;
      11'd894  : out_data_ref <= 8'h4a;
      11'd895  : out_data_ref <= 8'h6c;
      11'd896  : out_data_ref <= 8'hea;
      11'd897  : out_data_ref <= 8'ha6;
      11'd898  : out_data_ref <= 8'h5e;
      11'd899  : out_data_ref <= 8'h56;
      11'd900  : out_data_ref <= 8'h66;
      11'd901  : out_data_ref <= 8'h23;
      11'd902  : out_data_ref <= 8'h0a;
      11'd903  : out_data_ref <= 8'ha7;
      11'd904  : out_data_ref <= 8'h20;
      11'd905  : out_data_ref <= 8'h6a;
      11'd906  : out_data_ref <= 8'he7;
      11'd907  : out_data_ref <= 8'h8e;
      11'd908  : out_data_ref <= 8'hb1;
      11'd909  : out_data_ref <= 8'hb9;
      11'd910  : out_data_ref <= 8'h8c;
      11'd911  : out_data_ref <= 8'hb5;
      11'd912  : out_data_ref <= 8'h23;
      11'd913  : out_data_ref <= 8'h65;
      11'd914  : out_data_ref <= 8'h08;
      11'd915  : out_data_ref <= 8'he6;
      11'd916  : out_data_ref <= 8'h35;
      11'd917  : out_data_ref <= 8'h7e;
      11'd918  : out_data_ref <= 8'h18;
      11'd919  : out_data_ref <= 8'hcc;
      11'd920  : out_data_ref <= 8'hcf;
      11'd921  : out_data_ref <= 8'hae;
      11'd922  : out_data_ref <= 8'hc5;
      11'd923  : out_data_ref <= 8'h69;
      11'd924  : out_data_ref <= 8'h35;
      11'd925  : out_data_ref <= 8'h32;
      11'd926  : out_data_ref <= 8'hbe;
      11'd927  : out_data_ref <= 8'h4e;
      11'd928  : out_data_ref <= 8'he3;
      11'd929  : out_data_ref <= 8'h80;
      11'd930  : out_data_ref <= 8'h22;
      11'd931  : out_data_ref <= 8'hc4;
      11'd932  : out_data_ref <= 8'h8f;
      11'd933  : out_data_ref <= 8'he9;
      11'd934  : out_data_ref <= 8'h4f;
      11'd935  : out_data_ref <= 8'h62;
      11'd936  : out_data_ref <= 8'hb0;
      11'd937  : out_data_ref <= 8'h29;
      11'd938  : out_data_ref <= 8'h3a;
      11'd939  : out_data_ref <= 8'h08;
      11'd940  : out_data_ref <= 8'h8b;
      11'd941  : out_data_ref <= 8'hf4;
      11'd942  : out_data_ref <= 8'hd7;
      11'd943  : out_data_ref <= 8'h37;
      11'd944  : out_data_ref <= 8'hf4;
      11'd945  : out_data_ref <= 8'h87;
      11'd946  : out_data_ref <= 8'h48;
      11'd947  : out_data_ref <= 8'hf2;
      11'd948  : out_data_ref <= 8'h3b;
      11'd949  : out_data_ref <= 8'hcb;
      11'd950  : out_data_ref <= 8'h33;
      11'd951  : out_data_ref <= 8'h8b;
      11'd952  : out_data_ref <= 8'h58;
      11'd953  : out_data_ref <= 8'hb4;
      11'd954  : out_data_ref <= 8'hd6;
      11'd955  : out_data_ref <= 8'h66;
      11'd956  : out_data_ref <= 8'had;
      11'd957  : out_data_ref <= 8'h3c;
      11'd958  : out_data_ref <= 8'h64;
      11'd959  : out_data_ref <= 8'he9;
      11'd960  : out_data_ref <= 8'hec;
      11'd961  : out_data_ref <= 8'hd0;
      11'd962  : out_data_ref <= 8'h72;
      11'd963  : out_data_ref <= 8'h65;
      11'd964  : out_data_ref <= 8'hf9;
      11'd965  : out_data_ref <= 8'h71;
      11'd966  : out_data_ref <= 8'hb0;
      11'd967  : out_data_ref <= 8'h7a;
      11'd968  : out_data_ref <= 8'hf7;
      11'd969  : out_data_ref <= 8'h16;
      11'd970  : out_data_ref <= 8'hd4;
      11'd971  : out_data_ref <= 8'ha5;
      11'd972  : out_data_ref <= 8'hb7;
      11'd973  : out_data_ref <= 8'h19;
      11'd974  : out_data_ref <= 8'hc3;
      11'd975  : out_data_ref <= 8'hf5;
      11'd976  : out_data_ref <= 8'hfe;
      11'd977  : out_data_ref <= 8'h35;
      11'd978  : out_data_ref <= 8'h74;
      11'd979  : out_data_ref <= 8'h47;
      11'd980  : out_data_ref <= 8'h34;
      11'd981  : out_data_ref <= 8'hcb;
      11'd982  : out_data_ref <= 8'ha5;
      11'd983  : out_data_ref <= 8'h43;
      11'd984  : out_data_ref <= 8'h03;
      11'd985  : out_data_ref <= 8'h81;
      11'd986  : out_data_ref <= 8'h66;
      11'd987  : out_data_ref <= 8'h1e;
      11'd988  : out_data_ref <= 8'h37;
      11'd989  : out_data_ref <= 8'h2b;
      11'd990  : out_data_ref <= 8'h6f;
      11'd991  : out_data_ref <= 8'h65;
      11'd992  : out_data_ref <= 8'h10;
      11'd993  : out_data_ref <= 8'hd6;
      11'd994  : out_data_ref <= 8'h1b;
      11'd995  : out_data_ref <= 8'h11;
      11'd996  : out_data_ref <= 8'he4;
      11'd997  : out_data_ref <= 8'h69;
      11'd998  : out_data_ref <= 8'h7a;
      11'd999  : out_data_ref <= 8'h1a;
      11'd1000 : out_data_ref <= 8'h96;
      11'd1001 : out_data_ref <= 8'h15;
      11'd1002 : out_data_ref <= 8'h89;
      11'd1003 : out_data_ref <= 8'h94;
      11'd1004 : out_data_ref <= 8'h9d;
      11'd1005 : out_data_ref <= 8'hba;
      11'd1006 : out_data_ref <= 8'h53;
      11'd1007 : out_data_ref <= 8'hb5;
      11'd1008 : out_data_ref <= 8'hbc;
      11'd1009 : out_data_ref <= 8'h5b;
      11'd1010 : out_data_ref <= 8'hdb;
      11'd1011 : out_data_ref <= 8'h76;
      11'd1012 : out_data_ref <= 8'hfa;
      11'd1013 : out_data_ref <= 8'h09;
      11'd1014 : out_data_ref <= 8'h32;
      11'd1015 : out_data_ref <= 8'h43;
      11'd1016 : out_data_ref <= 8'h87;
      11'd1017 : out_data_ref <= 8'hd7;
      11'd1018 : out_data_ref <= 8'h99;
      11'd1019 : out_data_ref <= 8'h53;
      11'd1020 : out_data_ref <= 8'h65;
      11'd1021 : out_data_ref <= 8'h06;
      11'd1022 : out_data_ref <= 8'h18;
      11'd1023 : out_data_ref <= 8'h2e;
      11'd1024 : out_data_ref <= 8'hff;
      11'd1025 : out_data_ref <= 8'h70;
      11'd1026 : out_data_ref <= 8'h78;
      11'd1027 : out_data_ref <= 8'h03;
      11'd1028 : out_data_ref <= 8'h4b;
      11'd1029 : out_data_ref <= 8'h34;
      11'd1030 : out_data_ref <= 8'he1;
      11'd1031 : out_data_ref <= 8'hdd;
      11'd1032 : out_data_ref <= 8'hd2;
      11'd1033 : out_data_ref <= 8'h61;
      11'd1034 : out_data_ref <= 8'h2b;
      11'd1035 : out_data_ref <= 8'h0a;
      11'd1036 : out_data_ref <= 8'h40;
      11'd1037 : out_data_ref <= 8'he7;
      11'd1038 : out_data_ref <= 8'hf1;
      11'd1039 : out_data_ref <= 8'ha2;
      11'd1040 : out_data_ref <= 8'h94;
      11'd1041 : out_data_ref <= 8'hfb;
      11'd1042 : out_data_ref <= 8'ha8;
      11'd1043 : out_data_ref <= 8'h69;
      11'd1044 : out_data_ref <= 8'hda;
      11'd1045 : out_data_ref <= 8'h2e;
      11'd1046 : out_data_ref <= 8'h46;
      11'd1047 : out_data_ref <= 8'hc4;
      11'd1048 : out_data_ref <= 8'hc3;
      11'd1049 : out_data_ref <= 8'h6b;
      11'd1050 : out_data_ref <= 8'hb0;
      11'd1051 : out_data_ref <= 8'h8c;
      11'd1052 : out_data_ref <= 8'h7e;
      11'd1053 : out_data_ref <= 8'h9b;
      11'd1054 : out_data_ref <= 8'hef;
      11'd1055 : out_data_ref <= 8'h09;
      11'd1056 : out_data_ref <= 8'ha9;
      11'd1057 : out_data_ref <= 8'h44;
      11'd1058 : out_data_ref <= 8'h59;
      11'd1059 : out_data_ref <= 8'he8;
      11'd1060 : out_data_ref <= 8'hfc;
      11'd1061 : out_data_ref <= 8'h2d;
      11'd1062 : out_data_ref <= 8'h3c;
      11'd1063 : out_data_ref <= 8'hc5;
      11'd1064 : out_data_ref <= 8'h79;
      11'd1065 : out_data_ref <= 8'hd1;
      11'd1066 : out_data_ref <= 8'h52;
      11'd1067 : out_data_ref <= 8'h84;
      11'd1068 : out_data_ref <= 8'hdf;
      11'd1069 : out_data_ref <= 8'h1f;
      11'd1070 : out_data_ref <= 8'h19;
      11'd1071 : out_data_ref <= 8'hef;
      11'd1072 : out_data_ref <= 8'h77;
      11'd1073 : out_data_ref <= 8'he0;
      11'd1074 : out_data_ref <= 8'h30;
      11'd1075 : out_data_ref <= 8'h41;
      11'd1076 : out_data_ref <= 8'h51;
      11'd1077 : out_data_ref <= 8'h1a;
      11'd1078 : out_data_ref <= 8'hcc;
      11'd1079 : out_data_ref <= 8'h39;
      11'd1080 : out_data_ref <= 8'hbf;
      11'd1081 : out_data_ref <= 8'h9c;
      11'd1082 : out_data_ref <= 8'ha8;
      11'd1083 : out_data_ref <= 8'hac;
      11'd1084 : out_data_ref <= 8'h8d;
      11'd1085 : out_data_ref <= 8'he6;
      11'd1086 : out_data_ref <= 8'ha0;
      11'd1087 : out_data_ref <= 8'he5;
      11'd1088 : out_data_ref <= 8'hee;
      11'd1089 : out_data_ref <= 8'ha0;
      11'd1090 : out_data_ref <= 8'hbb;
      11'd1091 : out_data_ref <= 8'hd4;
      11'd1092 : out_data_ref <= 8'h28;
      11'd1093 : out_data_ref <= 8'h9b;
      11'd1094 : out_data_ref <= 8'h6d;
      11'd1095 : out_data_ref <= 8'hae;
      11'd1096 : out_data_ref <= 8'h38;
      11'd1097 : out_data_ref <= 8'he9;
      11'd1098 : out_data_ref <= 8'he8;
      11'd1099 : out_data_ref <= 8'h2e;
      11'd1100 : out_data_ref <= 8'hb5;
      11'd1101 : out_data_ref <= 8'h0a;
      11'd1102 : out_data_ref <= 8'h03;
      11'd1103 : out_data_ref <= 8'h97;
      11'd1104 : out_data_ref <= 8'hb3;
      11'd1105 : out_data_ref <= 8'hee;
      11'd1106 : out_data_ref <= 8'h6c;
      11'd1107 : out_data_ref <= 8'h52;
      11'd1108 : out_data_ref <= 8'hfb;
      11'd1109 : out_data_ref <= 8'hdc;
      11'd1110 : out_data_ref <= 8'h7d;
      11'd1111 : out_data_ref <= 8'hee;
      11'd1112 : out_data_ref <= 8'ha2;
      11'd1113 : out_data_ref <= 8'hc3;
      11'd1114 : out_data_ref <= 8'h76;
      11'd1115 : out_data_ref <= 8'h82;
      11'd1116 : out_data_ref <= 8'h5e;
      11'd1117 : out_data_ref <= 8'h89;
      11'd1118 : out_data_ref <= 8'h01;
      11'd1119 : out_data_ref <= 8'h6c;
      11'd1120 : out_data_ref <= 8'h85;
      11'd1121 : out_data_ref <= 8'h9b;
      11'd1122 : out_data_ref <= 8'h09;
      11'd1123 : out_data_ref <= 8'h48;
      11'd1124 : out_data_ref <= 8'h85;
      11'd1125 : out_data_ref <= 8'h48;
      11'd1126 : out_data_ref <= 8'hbf;
      11'd1127 : out_data_ref <= 8'h76;
      11'd1128 : out_data_ref <= 8'hca;
      11'd1129 : out_data_ref <= 8'h62;
      11'd1130 : out_data_ref <= 8'hd6;
      11'd1131 : out_data_ref <= 8'h96;
      11'd1132 : out_data_ref <= 8'hdf;
      11'd1133 : out_data_ref <= 8'h94;
      11'd1134 : out_data_ref <= 8'ha6;
      11'd1135 : out_data_ref <= 8'h1e;
      11'd1136 : out_data_ref <= 8'h8f;
      11'd1137 : out_data_ref <= 8'h0e;
      11'd1138 : out_data_ref <= 8'h13;
      11'd1139 : out_data_ref <= 8'hc6;
      11'd1140 : out_data_ref <= 8'h9e;
      11'd1141 : out_data_ref <= 8'he8;
      11'd1142 : out_data_ref <= 8'h16;
      11'd1143 : out_data_ref <= 8'hce;
      11'd1144 : out_data_ref <= 8'h5a;
      11'd1145 : out_data_ref <= 8'ha2;
      11'd1146 : out_data_ref <= 8'h76;
      11'd1147 : out_data_ref <= 8'h89;
      11'd1148 : out_data_ref <= 8'h87;
      11'd1149 : out_data_ref <= 8'hb0;
      11'd1150 : out_data_ref <= 8'ha7;
      11'd1151 : out_data_ref <= 8'h82;
      11'd1152 : out_data_ref <= 8'hd7;
      11'd1153 : out_data_ref <= 8'h4c;
      11'd1154 : out_data_ref <= 8'h67;
      11'd1155 : out_data_ref <= 8'h3e;
      11'd1156 : out_data_ref <= 8'hc0;
      11'd1157 : out_data_ref <= 8'h05;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
