module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam R_LEN = 'd1013;
  localparam R_DEPTH = 'd10;
  localparam B_LEN = 'd1623;
  localparam B_DEPTH = 'd11;

  input              clk;
  input      [ 9: 0] in_addr;
  output reg [13: 0] in_data;
  input      [10: 0] out_addr;
  output reg [ 7: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      10'd0    : in_data <= 14'h1699; // 'd5785
      10'd1    : in_data <= 14'h169f; // 'd5791
      10'd2    : in_data <= 14'h1b32; // 'd6962
      10'd3    : in_data <= 14'h176a; // 'd5994
      10'd4    : in_data <= 14'h1391; // 'd5009
      10'd5    : in_data <= 14'h0be8; // 'd3048
      10'd6    : in_data <= 14'h1233; // 'd4659
      10'd7    : in_data <= 14'h03ad; // 'd941
      10'd8    : in_data <= 14'h054a; // 'd1354
      10'd9    : in_data <= 14'h0844; // 'd2116
      10'd10   : in_data <= 14'h142a; // 'd5162
      10'd11   : in_data <= 14'h12d3; // 'd4819
      10'd12   : in_data <= 14'h1939; // 'd6457
      10'd13   : in_data <= 14'h12d2; // 'd4818
      10'd14   : in_data <= 14'h1b58; // 'd7000
      10'd15   : in_data <= 14'h0ae0; // 'd2784
      10'd16   : in_data <= 14'h18a5; // 'd6309
      10'd17   : in_data <= 14'h0496; // 'd1174
      10'd18   : in_data <= 14'h151a; // 'd5402
      10'd19   : in_data <= 14'h0fde; // 'd4062
      10'd20   : in_data <= 14'h0ab2; // 'd2738
      10'd21   : in_data <= 14'h0d23; // 'd3363
      10'd22   : in_data <= 14'h0bb3; // 'd2995
      10'd23   : in_data <= 14'h035a; // 'd858
      10'd24   : in_data <= 14'h111c; // 'd4380
      10'd25   : in_data <= 14'h039e; // 'd926
      10'd26   : in_data <= 14'h0cd4; // 'd3284
      10'd27   : in_data <= 14'h1b80; // 'd7040
      10'd28   : in_data <= 14'h0fea; // 'd4074
      10'd29   : in_data <= 14'h0750; // 'd1872
      10'd30   : in_data <= 14'h1379; // 'd4985
      10'd31   : in_data <= 14'h0ebe; // 'd3774
      10'd32   : in_data <= 14'h0c32; // 'd3122
      10'd33   : in_data <= 14'h16d2; // 'd5842
      10'd34   : in_data <= 14'h0022; // 'd34
      10'd35   : in_data <= 14'h0834; // 'd2100
      10'd36   : in_data <= 14'h0cbd; // 'd3261
      10'd37   : in_data <= 14'h0afc; // 'd2812
      10'd38   : in_data <= 14'h0e40; // 'd3648
      10'd39   : in_data <= 14'h01ee; // 'd494
      10'd40   : in_data <= 14'h12b0; // 'd4784
      10'd41   : in_data <= 14'h1b52; // 'd6994
      10'd42   : in_data <= 14'h13cd; // 'd5069
      10'd43   : in_data <= 14'h038b; // 'd907
      10'd44   : in_data <= 14'h0a49; // 'd2633
      10'd45   : in_data <= 14'h1445; // 'd5189
      10'd46   : in_data <= 14'h1452; // 'd5202
      10'd47   : in_data <= 14'h12dd; // 'd4829
      10'd48   : in_data <= 14'h186a; // 'd6250
      10'd49   : in_data <= 14'h0eee; // 'd3822
      10'd50   : in_data <= 14'h0fa0; // 'd4000
      10'd51   : in_data <= 14'h0b10; // 'd2832
      10'd52   : in_data <= 14'h0e4f; // 'd3663
      10'd53   : in_data <= 14'h0965; // 'd2405
      10'd54   : in_data <= 14'h0838; // 'd2104
      10'd55   : in_data <= 14'h11f5; // 'd4597
      10'd56   : in_data <= 14'h0d0f; // 'd3343
      10'd57   : in_data <= 14'h0312; // 'd786
      10'd58   : in_data <= 14'h08db; // 'd2267
      10'd59   : in_data <= 14'h049a; // 'd1178
      10'd60   : in_data <= 14'h054b; // 'd1355
      10'd61   : in_data <= 14'h1249; // 'd4681
      10'd62   : in_data <= 14'h1100; // 'd4352
      10'd63   : in_data <= 14'h165d; // 'd5725
      10'd64   : in_data <= 14'h08f9; // 'd2297
      10'd65   : in_data <= 14'h0d63; // 'd3427
      10'd66   : in_data <= 14'h0e07; // 'd3591
      10'd67   : in_data <= 14'h12ea; // 'd4842
      10'd68   : in_data <= 14'h1b90; // 'd7056
      10'd69   : in_data <= 14'h1a1e; // 'd6686
      10'd70   : in_data <= 14'h0bd2; // 'd3026
      10'd71   : in_data <= 14'h1396; // 'd5014
      10'd72   : in_data <= 14'h1aed; // 'd6893
      10'd73   : in_data <= 14'h12a8; // 'd4776
      10'd74   : in_data <= 14'h0a61; // 'd2657
      10'd75   : in_data <= 14'h184a; // 'd6218
      10'd76   : in_data <= 14'h1516; // 'd5398
      10'd77   : in_data <= 14'h0021; // 'd33
      10'd78   : in_data <= 14'h01fa; // 'd506
      10'd79   : in_data <= 14'h0984; // 'd2436
      10'd80   : in_data <= 14'h0957; // 'd2391
      10'd81   : in_data <= 14'h1077; // 'd4215
      10'd82   : in_data <= 14'h051f; // 'd1311
      10'd83   : in_data <= 14'h1029; // 'd4137
      10'd84   : in_data <= 14'h0a6e; // 'd2670
      10'd85   : in_data <= 14'h0b5c; // 'd2908
      10'd86   : in_data <= 14'h19d8; // 'd6616
      10'd87   : in_data <= 14'h1395; // 'd5013
      10'd88   : in_data <= 14'h0f32; // 'd3890
      10'd89   : in_data <= 14'h0402; // 'd1026
      10'd90   : in_data <= 14'h1233; // 'd4659
      10'd91   : in_data <= 14'h09fb; // 'd2555
      10'd92   : in_data <= 14'h12bd; // 'd4797
      10'd93   : in_data <= 14'h1020; // 'd4128
      10'd94   : in_data <= 14'h08ac; // 'd2220
      10'd95   : in_data <= 14'h1837; // 'd6199
      10'd96   : in_data <= 14'h006a; // 'd106
      10'd97   : in_data <= 14'h109a; // 'd4250
      10'd98   : in_data <= 14'h0e25; // 'd3621
      10'd99   : in_data <= 14'h19fe; // 'd6654
      10'd100  : in_data <= 14'h1803; // 'd6147
      10'd101  : in_data <= 14'h19c0; // 'd6592
      10'd102  : in_data <= 14'h0165; // 'd357
      10'd103  : in_data <= 14'h1133; // 'd4403
      10'd104  : in_data <= 14'h0688; // 'd1672
      10'd105  : in_data <= 14'h1683; // 'd5763
      10'd106  : in_data <= 14'h035e; // 'd862
      10'd107  : in_data <= 14'h06d8; // 'd1752
      10'd108  : in_data <= 14'h1b22; // 'd6946
      10'd109  : in_data <= 14'h0587; // 'd1415
      10'd110  : in_data <= 14'h177c; // 'd6012
      10'd111  : in_data <= 14'h103e; // 'd4158
      10'd112  : in_data <= 14'h029c; // 'd668
      10'd113  : in_data <= 14'h0777; // 'd1911
      10'd114  : in_data <= 14'h198a; // 'd6538
      10'd115  : in_data <= 14'h17c1; // 'd6081
      10'd116  : in_data <= 14'h123f; // 'd4671
      10'd117  : in_data <= 14'h02c9; // 'd713
      10'd118  : in_data <= 14'h06b7; // 'd1719
      10'd119  : in_data <= 14'h145a; // 'd5210
      10'd120  : in_data <= 14'h030e; // 'd782
      10'd121  : in_data <= 14'h08ea; // 'd2282
      10'd122  : in_data <= 14'h0475; // 'd1141
      10'd123  : in_data <= 14'h119c; // 'd4508
      10'd124  : in_data <= 14'h06f2; // 'd1778
      10'd125  : in_data <= 14'h0514; // 'd1300
      10'd126  : in_data <= 14'h0096; // 'd150
      10'd127  : in_data <= 14'h1540; // 'd5440
      10'd128  : in_data <= 14'h119a; // 'd4506
      10'd129  : in_data <= 14'h1905; // 'd6405
      10'd130  : in_data <= 14'h164a; // 'd5706
      10'd131  : in_data <= 14'h0c22; // 'd3106
      10'd132  : in_data <= 14'h08ef; // 'd2287
      10'd133  : in_data <= 14'h0f8e; // 'd3982
      10'd134  : in_data <= 14'h070f; // 'd1807
      10'd135  : in_data <= 14'h1501; // 'd5377
      10'd136  : in_data <= 14'h0cf2; // 'd3314
      10'd137  : in_data <= 14'h0cc6; // 'd3270
      10'd138  : in_data <= 14'h17a2; // 'd6050
      10'd139  : in_data <= 14'h0eb6; // 'd3766
      10'd140  : in_data <= 14'h0abb; // 'd2747
      10'd141  : in_data <= 14'h13af; // 'd5039
      10'd142  : in_data <= 14'h14ac; // 'd5292
      10'd143  : in_data <= 14'h0851; // 'd2129
      10'd144  : in_data <= 14'h17f1; // 'd6129
      10'd145  : in_data <= 14'h10d0; // 'd4304
      10'd146  : in_data <= 14'h1831; // 'd6193
      10'd147  : in_data <= 14'h01c2; // 'd450
      10'd148  : in_data <= 14'h1a67; // 'd6759
      10'd149  : in_data <= 14'h1156; // 'd4438
      10'd150  : in_data <= 14'h1323; // 'd4899
      10'd151  : in_data <= 14'h06a7; // 'd1703
      10'd152  : in_data <= 14'h0fca; // 'd4042
      10'd153  : in_data <= 14'h0603; // 'd1539
      10'd154  : in_data <= 14'h1913; // 'd6419
      10'd155  : in_data <= 14'h19bd; // 'd6589
      10'd156  : in_data <= 14'h09d8; // 'd2520
      10'd157  : in_data <= 14'h188c; // 'd6284
      10'd158  : in_data <= 14'h0942; // 'd2370
      10'd159  : in_data <= 14'h178e; // 'd6030
      10'd160  : in_data <= 14'h03e5; // 'd997
      10'd161  : in_data <= 14'h14e0; // 'd5344
      10'd162  : in_data <= 14'h02ba; // 'd698
      10'd163  : in_data <= 14'h165b; // 'd5723
      10'd164  : in_data <= 14'h0f2a; // 'd3882
      10'd165  : in_data <= 14'h178d; // 'd6029
      10'd166  : in_data <= 14'h0947; // 'd2375
      10'd167  : in_data <= 14'h19e2; // 'd6626
      10'd168  : in_data <= 14'h0f7b; // 'd3963
      10'd169  : in_data <= 14'h038d; // 'd909
      10'd170  : in_data <= 14'h13a2; // 'd5026
      10'd171  : in_data <= 14'h0b51; // 'd2897
      10'd172  : in_data <= 14'h13a6; // 'd5030
      10'd173  : in_data <= 14'h03f3; // 'd1011
      10'd174  : in_data <= 14'h0c31; // 'd3121
      10'd175  : in_data <= 14'h0416; // 'd1046
      10'd176  : in_data <= 14'h06b8; // 'd1720
      10'd177  : in_data <= 14'h005f; // 'd95
      10'd178  : in_data <= 14'h0709; // 'd1801
      10'd179  : in_data <= 14'h0307; // 'd775
      10'd180  : in_data <= 14'h073b; // 'd1851
      10'd181  : in_data <= 14'h13d8; // 'd5080
      10'd182  : in_data <= 14'h101b; // 'd4123
      10'd183  : in_data <= 14'h095b; // 'd2395
      10'd184  : in_data <= 14'h1a4b; // 'd6731
      10'd185  : in_data <= 14'h1b5c; // 'd7004
      10'd186  : in_data <= 14'h1a5a; // 'd6746
      10'd187  : in_data <= 14'h068e; // 'd1678
      10'd188  : in_data <= 14'h0213; // 'd531
      10'd189  : in_data <= 14'h0f5d; // 'd3933
      10'd190  : in_data <= 14'h0ede; // 'd3806
      10'd191  : in_data <= 14'h163e; // 'd5694
      10'd192  : in_data <= 14'h0a18; // 'd2584
      10'd193  : in_data <= 14'h0204; // 'd516
      10'd194  : in_data <= 14'h0dd0; // 'd3536
      10'd195  : in_data <= 14'h167e; // 'd5758
      10'd196  : in_data <= 14'h0eb9; // 'd3769
      10'd197  : in_data <= 14'h01f6; // 'd502
      10'd198  : in_data <= 14'h0c73; // 'd3187
      10'd199  : in_data <= 14'h1239; // 'd4665
      10'd200  : in_data <= 14'h09e4; // 'd2532
      10'd201  : in_data <= 14'h11f5; // 'd4597
      10'd202  : in_data <= 14'h1b1b; // 'd6939
      10'd203  : in_data <= 14'h0294; // 'd660
      10'd204  : in_data <= 14'h177e; // 'd6014
      10'd205  : in_data <= 14'h0013; // 'd19
      10'd206  : in_data <= 14'h0b54; // 'd2900
      10'd207  : in_data <= 14'h114e; // 'd4430
      10'd208  : in_data <= 14'h0fe6; // 'd4070
      10'd209  : in_data <= 14'h1a05; // 'd6661
      10'd210  : in_data <= 14'h10a4; // 'd4260
      10'd211  : in_data <= 14'h1591; // 'd5521
      10'd212  : in_data <= 14'h0b15; // 'd2837
      10'd213  : in_data <= 14'h1595; // 'd5525
      10'd214  : in_data <= 14'h11fb; // 'd4603
      10'd215  : in_data <= 14'h004c; // 'd76
      10'd216  : in_data <= 14'h1521; // 'd5409
      10'd217  : in_data <= 14'h0a3e; // 'd2622
      10'd218  : in_data <= 14'h150d; // 'd5389
      10'd219  : in_data <= 14'h1517; // 'd5399
      10'd220  : in_data <= 14'h0405; // 'd1029
      10'd221  : in_data <= 14'h0e02; // 'd3586
      10'd222  : in_data <= 14'h157e; // 'd5502
      10'd223  : in_data <= 14'h0a47; // 'd2631
      10'd224  : in_data <= 14'h1866; // 'd6246
      10'd225  : in_data <= 14'h04a4; // 'd1188
      10'd226  : in_data <= 14'h1b02; // 'd6914
      10'd227  : in_data <= 14'h01d9; // 'd473
      10'd228  : in_data <= 14'h0cb4; // 'd3252
      10'd229  : in_data <= 14'h0220; // 'd544
      10'd230  : in_data <= 14'h0a6f; // 'd2671
      10'd231  : in_data <= 14'h13dc; // 'd5084
      10'd232  : in_data <= 14'h1784; // 'd6020
      10'd233  : in_data <= 14'h050d; // 'd1293
      10'd234  : in_data <= 14'h04bf; // 'd1215
      10'd235  : in_data <= 14'h03a1; // 'd929
      10'd236  : in_data <= 14'h1106; // 'd4358
      10'd237  : in_data <= 14'h003f; // 'd63
      10'd238  : in_data <= 14'h0c9d; // 'd3229
      10'd239  : in_data <= 14'h0434; // 'd1076
      10'd240  : in_data <= 14'h133f; // 'd4927
      10'd241  : in_data <= 14'h015d; // 'd349
      10'd242  : in_data <= 14'h0ff4; // 'd4084
      10'd243  : in_data <= 14'h18d2; // 'd6354
      10'd244  : in_data <= 14'h0048; // 'd72
      10'd245  : in_data <= 14'h01a5; // 'd421
      10'd246  : in_data <= 14'h0bdd; // 'd3037
      10'd247  : in_data <= 14'h17a6; // 'd6054
      10'd248  : in_data <= 14'h1ad7; // 'd6871
      10'd249  : in_data <= 14'h0b22; // 'd2850
      10'd250  : in_data <= 14'h11f4; // 'd4596
      10'd251  : in_data <= 14'h1919; // 'd6425
      10'd252  : in_data <= 14'h07d5; // 'd2005
      10'd253  : in_data <= 14'h07d4; // 'd2004
      10'd254  : in_data <= 14'h082e; // 'd2094
      10'd255  : in_data <= 14'h1118; // 'd4376
      10'd256  : in_data <= 14'h0354; // 'd852
      10'd257  : in_data <= 14'h0090; // 'd144
      10'd258  : in_data <= 14'h16d3; // 'd5843
      10'd259  : in_data <= 14'h07a5; // 'd1957
      10'd260  : in_data <= 14'h1add; // 'd6877
      10'd261  : in_data <= 14'h0bbf; // 'd3007
      10'd262  : in_data <= 14'h01e5; // 'd485
      10'd263  : in_data <= 14'h1aa2; // 'd6818
      10'd264  : in_data <= 14'h05b6; // 'd1462
      10'd265  : in_data <= 14'h0336; // 'd822
      10'd266  : in_data <= 14'h10bd; // 'd4285
      10'd267  : in_data <= 14'h1940; // 'd6464
      10'd268  : in_data <= 14'h1491; // 'd5265
      10'd269  : in_data <= 14'h1210; // 'd4624
      10'd270  : in_data <= 14'h13ba; // 'd5050
      10'd271  : in_data <= 14'h1973; // 'd6515
      10'd272  : in_data <= 14'h116a; // 'd4458
      10'd273  : in_data <= 14'h0f76; // 'd3958
      10'd274  : in_data <= 14'h151c; // 'd5404
      10'd275  : in_data <= 14'h18b9; // 'd6329
      10'd276  : in_data <= 14'h0036; // 'd54
      10'd277  : in_data <= 14'h132c; // 'd4908
      10'd278  : in_data <= 14'h0199; // 'd409
      10'd279  : in_data <= 14'h043e; // 'd1086
      10'd280  : in_data <= 14'h03f9; // 'd1017
      10'd281  : in_data <= 14'h0876; // 'd2166
      10'd282  : in_data <= 14'h15e6; // 'd5606
      10'd283  : in_data <= 14'h00e7; // 'd231
      10'd284  : in_data <= 14'h1518; // 'd5400
      10'd285  : in_data <= 14'h0142; // 'd322
      10'd286  : in_data <= 14'h1aad; // 'd6829
      10'd287  : in_data <= 14'h1252; // 'd4690
      10'd288  : in_data <= 14'h13b0; // 'd5040
      10'd289  : in_data <= 14'h1944; // 'd6468
      10'd290  : in_data <= 14'h07c3; // 'd1987
      10'd291  : in_data <= 14'h060c; // 'd1548
      10'd292  : in_data <= 14'h14db; // 'd5339
      10'd293  : in_data <= 14'h014b; // 'd331
      10'd294  : in_data <= 14'h0999; // 'd2457
      10'd295  : in_data <= 14'h13cf; // 'd5071
      10'd296  : in_data <= 14'h01f7; // 'd503
      10'd297  : in_data <= 14'h0ce1; // 'd3297
      10'd298  : in_data <= 14'h0250; // 'd592
      10'd299  : in_data <= 14'h11be; // 'd4542
      10'd300  : in_data <= 14'h0748; // 'd1864
      10'd301  : in_data <= 14'h1b50; // 'd6992
      10'd302  : in_data <= 14'h0b7b; // 'd2939
      10'd303  : in_data <= 14'h05b0; // 'd1456
      10'd304  : in_data <= 14'h0dee; // 'd3566
      10'd305  : in_data <= 14'h0c54; // 'd3156
      10'd306  : in_data <= 14'h07e4; // 'd2020
      10'd307  : in_data <= 14'h15a5; // 'd5541
      10'd308  : in_data <= 14'h0f98; // 'd3992
      10'd309  : in_data <= 14'h12c0; // 'd4800
      10'd310  : in_data <= 14'h0f79; // 'd3961
      10'd311  : in_data <= 14'h0942; // 'd2370
      10'd312  : in_data <= 14'h0121; // 'd289
      10'd313  : in_data <= 14'h09f1; // 'd2545
      10'd314  : in_data <= 14'h1607; // 'd5639
      10'd315  : in_data <= 14'h0207; // 'd519
      10'd316  : in_data <= 14'h0169; // 'd361
      10'd317  : in_data <= 14'h132a; // 'd4906
      10'd318  : in_data <= 14'h023d; // 'd573
      10'd319  : in_data <= 14'h0704; // 'd1796
      10'd320  : in_data <= 14'h105a; // 'd4186
      10'd321  : in_data <= 14'h02fc; // 'd764
      10'd322  : in_data <= 14'h1137; // 'd4407
      10'd323  : in_data <= 14'h08bf; // 'd2239
      10'd324  : in_data <= 14'h00a6; // 'd166
      10'd325  : in_data <= 14'h19a3; // 'd6563
      10'd326  : in_data <= 14'h02f0; // 'd752
      10'd327  : in_data <= 14'h1573; // 'd5491
      10'd328  : in_data <= 14'h158c; // 'd5516
      10'd329  : in_data <= 14'h17b2; // 'd6066
      10'd330  : in_data <= 14'h00bc; // 'd188
      10'd331  : in_data <= 14'h1ba8; // 'd7080
      10'd332  : in_data <= 14'h1521; // 'd5409
      10'd333  : in_data <= 14'h1992; // 'd6546
      10'd334  : in_data <= 14'h09e9; // 'd2537
      10'd335  : in_data <= 14'h05f7; // 'd1527
      10'd336  : in_data <= 14'h1b54; // 'd6996
      10'd337  : in_data <= 14'h1a8d; // 'd6797
      10'd338  : in_data <= 14'h06ea; // 'd1770
      10'd339  : in_data <= 14'h0d21; // 'd3361
      10'd340  : in_data <= 14'h118a; // 'd4490
      10'd341  : in_data <= 14'h1327; // 'd4903
      10'd342  : in_data <= 14'h084a; // 'd2122
      10'd343  : in_data <= 14'h0af3; // 'd2803
      10'd344  : in_data <= 14'h1832; // 'd6194
      10'd345  : in_data <= 14'h0ef9; // 'd3833
      10'd346  : in_data <= 14'h0646; // 'd1606
      10'd347  : in_data <= 14'h18da; // 'd6362
      10'd348  : in_data <= 14'h03fc; // 'd1020
      10'd349  : in_data <= 14'h02dc; // 'd732
      10'd350  : in_data <= 14'h02c0; // 'd704
      10'd351  : in_data <= 14'h07b3; // 'd1971
      10'd352  : in_data <= 14'h1834; // 'd6196
      10'd353  : in_data <= 14'h1b81; // 'd7041
      10'd354  : in_data <= 14'h0ca7; // 'd3239
      10'd355  : in_data <= 14'h0491; // 'd1169
      10'd356  : in_data <= 14'h11e0; // 'd4576
      10'd357  : in_data <= 14'h13d4; // 'd5076
      10'd358  : in_data <= 14'h0241; // 'd577
      10'd359  : in_data <= 14'h0030; // 'd48
      10'd360  : in_data <= 14'h1324; // 'd4900
      10'd361  : in_data <= 14'h0064; // 'd100
      10'd362  : in_data <= 14'h046c; // 'd1132
      10'd363  : in_data <= 14'h18de; // 'd6366
      10'd364  : in_data <= 14'h08e4; // 'd2276
      10'd365  : in_data <= 14'h148a; // 'd5258
      10'd366  : in_data <= 14'h19e5; // 'd6629
      10'd367  : in_data <= 14'h0235; // 'd565
      10'd368  : in_data <= 14'h0354; // 'd852
      10'd369  : in_data <= 14'h1511; // 'd5393
      10'd370  : in_data <= 14'h1b67; // 'd7015
      10'd371  : in_data <= 14'h0bd1; // 'd3025
      10'd372  : in_data <= 14'h02e4; // 'd740
      10'd373  : in_data <= 14'h0ad9; // 'd2777
      10'd374  : in_data <= 14'h0cb7; // 'd3255
      10'd375  : in_data <= 14'h0488; // 'd1160
      10'd376  : in_data <= 14'h0a8d; // 'd2701
      10'd377  : in_data <= 14'h18e6; // 'd6374
      10'd378  : in_data <= 14'h0fad; // 'd4013
      10'd379  : in_data <= 14'h08fc; // 'd2300
      10'd380  : in_data <= 14'h03d6; // 'd982
      10'd381  : in_data <= 14'h0ef5; // 'd3829
      10'd382  : in_data <= 14'h00a3; // 'd163
      10'd383  : in_data <= 14'h0ed5; // 'd3797
      10'd384  : in_data <= 14'h086a; // 'd2154
      10'd385  : in_data <= 14'h0f45; // 'd3909
      10'd386  : in_data <= 14'h0135; // 'd309
      10'd387  : in_data <= 14'h1701; // 'd5889
      10'd388  : in_data <= 14'h0d8e; // 'd3470
      10'd389  : in_data <= 14'h0488; // 'd1160
      10'd390  : in_data <= 14'h0ab5; // 'd2741
      10'd391  : in_data <= 14'h18c2; // 'd6338
      10'd392  : in_data <= 14'h05d1; // 'd1489
      10'd393  : in_data <= 14'h095c; // 'd2396
      10'd394  : in_data <= 14'h167c; // 'd5756
      10'd395  : in_data <= 14'h09a6; // 'd2470
      10'd396  : in_data <= 14'h125f; // 'd4703
      10'd397  : in_data <= 14'h070e; // 'd1806
      10'd398  : in_data <= 14'h0c82; // 'd3202
      10'd399  : in_data <= 14'h1983; // 'd6531
      10'd400  : in_data <= 14'h092f; // 'd2351
      10'd401  : in_data <= 14'h07b0; // 'd1968
      10'd402  : in_data <= 14'h02f7; // 'd759
      10'd403  : in_data <= 14'h0e95; // 'd3733
      10'd404  : in_data <= 14'h057d; // 'd1405
      10'd405  : in_data <= 14'h1160; // 'd4448
      10'd406  : in_data <= 14'h0363; // 'd867
      10'd407  : in_data <= 14'h0799; // 'd1945
      10'd408  : in_data <= 14'h18c3; // 'd6339
      10'd409  : in_data <= 14'h0352; // 'd850
      10'd410  : in_data <= 14'h0549; // 'd1353
      10'd411  : in_data <= 14'h0b2a; // 'd2858
      10'd412  : in_data <= 14'h0c2e; // 'd3118
      10'd413  : in_data <= 14'h0b1d; // 'd2845
      10'd414  : in_data <= 14'h119d; // 'd4509
      10'd415  : in_data <= 14'h05b9; // 'd1465
      10'd416  : in_data <= 14'h0db1; // 'd3505
      10'd417  : in_data <= 14'h0360; // 'd864
      10'd418  : in_data <= 14'h1bc9; // 'd7113
      10'd419  : in_data <= 14'h108b; // 'd4235
      10'd420  : in_data <= 14'h1099; // 'd4249
      10'd421  : in_data <= 14'h0abc; // 'd2748
      10'd422  : in_data <= 14'h0079; // 'd121
      10'd423  : in_data <= 14'h136a; // 'd4970
      10'd424  : in_data <= 14'h0035; // 'd53
      10'd425  : in_data <= 14'h0b47; // 'd2887
      10'd426  : in_data <= 14'h11d1; // 'd4561
      10'd427  : in_data <= 14'h0328; // 'd808
      10'd428  : in_data <= 14'h053b; // 'd1339
      10'd429  : in_data <= 14'h1924; // 'd6436
      10'd430  : in_data <= 14'h0ea2; // 'd3746
      10'd431  : in_data <= 14'h0f61; // 'd3937
      10'd432  : in_data <= 14'h1425; // 'd5157
      10'd433  : in_data <= 14'h0b97; // 'd2967
      10'd434  : in_data <= 14'h1412; // 'd5138
      10'd435  : in_data <= 14'h1864; // 'd6244
      10'd436  : in_data <= 14'h1591; // 'd5521
      10'd437  : in_data <= 14'h1289; // 'd4745
      10'd438  : in_data <= 14'h1b52; // 'd6994
      10'd439  : in_data <= 14'h19d3; // 'd6611
      10'd440  : in_data <= 14'h0537; // 'd1335
      10'd441  : in_data <= 14'h0148; // 'd328
      10'd442  : in_data <= 14'h052c; // 'd1324
      10'd443  : in_data <= 14'h0ef4; // 'd3828
      10'd444  : in_data <= 14'h02ee; // 'd750
      10'd445  : in_data <= 14'h1514; // 'd5396
      10'd446  : in_data <= 14'h062a; // 'd1578
      10'd447  : in_data <= 14'h1054; // 'd4180
      10'd448  : in_data <= 14'h159c; // 'd5532
      10'd449  : in_data <= 14'h0cf3; // 'd3315
      10'd450  : in_data <= 14'h186c; // 'd6252
      10'd451  : in_data <= 14'h1031; // 'd4145
      10'd452  : in_data <= 14'h0ae4; // 'd2788
      10'd453  : in_data <= 14'h0653; // 'd1619
      10'd454  : in_data <= 14'h0be5; // 'd3045
      10'd455  : in_data <= 14'h099a; // 'd2458
      10'd456  : in_data <= 14'h0eb5; // 'd3765
      10'd457  : in_data <= 14'h17ac; // 'd6060
      10'd458  : in_data <= 14'h07de; // 'd2014
      10'd459  : in_data <= 14'h1715; // 'd5909
      10'd460  : in_data <= 14'h157a; // 'd5498
      10'd461  : in_data <= 14'h0837; // 'd2103
      10'd462  : in_data <= 14'h1a16; // 'd6678
      10'd463  : in_data <= 14'h05c2; // 'd1474
      10'd464  : in_data <= 14'h078a; // 'd1930
      10'd465  : in_data <= 14'h0d22; // 'd3362
      10'd466  : in_data <= 14'h1a3f; // 'd6719
      10'd467  : in_data <= 14'h0ab7; // 'd2743
      10'd468  : in_data <= 14'h0d9e; // 'd3486
      10'd469  : in_data <= 14'h0f24; // 'd3876
      10'd470  : in_data <= 14'h0d2a; // 'd3370
      10'd471  : in_data <= 14'h0d16; // 'd3350
      10'd472  : in_data <= 14'h0704; // 'd1796
      10'd473  : in_data <= 14'h0f04; // 'd3844
      10'd474  : in_data <= 14'h1b69; // 'd7017
      10'd475  : in_data <= 14'h00eb; // 'd235
      10'd476  : in_data <= 14'h0c52; // 'd3154
      10'd477  : in_data <= 14'h0daf; // 'd3503
      10'd478  : in_data <= 14'h0a6b; // 'd2667
      10'd479  : in_data <= 14'h09bf; // 'd2495
      10'd480  : in_data <= 14'h06e5; // 'd1765
      10'd481  : in_data <= 14'h182a; // 'd6186
      10'd482  : in_data <= 14'h0209; // 'd521
      10'd483  : in_data <= 14'h17c7; // 'd6087
      10'd484  : in_data <= 14'h1af2; // 'd6898
      10'd485  : in_data <= 14'h0d9d; // 'd3485
      10'd486  : in_data <= 14'h0ba4; // 'd2980
      10'd487  : in_data <= 14'h1bcf; // 'd7119
      10'd488  : in_data <= 14'h07b4; // 'd1972
      10'd489  : in_data <= 14'h168e; // 'd5774
      10'd490  : in_data <= 14'h15a7; // 'd5543
      10'd491  : in_data <= 14'h156e; // 'd5486
      10'd492  : in_data <= 14'h0d9d; // 'd3485
      10'd493  : in_data <= 14'h0108; // 'd264
      10'd494  : in_data <= 14'h141b; // 'd5147
      10'd495  : in_data <= 14'h06dc; // 'd1756
      10'd496  : in_data <= 14'h0c63; // 'd3171
      10'd497  : in_data <= 14'h050e; // 'd1294
      10'd498  : in_data <= 14'h1b08; // 'd6920
      10'd499  : in_data <= 14'h01d7; // 'd471
      10'd500  : in_data <= 14'h1a46; // 'd6726
      10'd501  : in_data <= 14'h068b; // 'd1675
      10'd502  : in_data <= 14'h0b72; // 'd2930
      10'd503  : in_data <= 14'h0457; // 'd1111
      10'd504  : in_data <= 14'h054b; // 'd1355
      10'd505  : in_data <= 14'h1b95; // 'd7061
      10'd506  : in_data <= 14'h04e0; // 'd1248
      10'd507  : in_data <= 14'h19c3; // 'd6595
      10'd508  : in_data <= 14'h0336; // 'd822
      10'd509  : in_data <= 14'h01e9; // 'd489
      10'd510  : in_data <= 14'h0dfd; // 'd3581
      10'd511  : in_data <= 14'h1478; // 'd5240
      10'd512  : in_data <= 14'h093e; // 'd2366
      10'd513  : in_data <= 14'h0974; // 'd2420
      10'd514  : in_data <= 14'h1499; // 'd5273
      10'd515  : in_data <= 14'h0ef0; // 'd3824
      10'd516  : in_data <= 14'h058c; // 'd1420
      10'd517  : in_data <= 14'h101d; // 'd4125
      10'd518  : in_data <= 14'h128c; // 'd4748
      10'd519  : in_data <= 14'h1728; // 'd5928
      10'd520  : in_data <= 14'h18ce; // 'd6350
      10'd521  : in_data <= 14'h1884; // 'd6276
      10'd522  : in_data <= 14'h1561; // 'd5473
      10'd523  : in_data <= 14'h01e7; // 'd487
      10'd524  : in_data <= 14'h0aa2; // 'd2722
      10'd525  : in_data <= 14'h13d7; // 'd5079
      10'd526  : in_data <= 14'h18c5; // 'd6341
      10'd527  : in_data <= 14'h17f2; // 'd6130
      10'd528  : in_data <= 14'h1267; // 'd4711
      10'd529  : in_data <= 14'h01e5; // 'd485
      10'd530  : in_data <= 14'h1895; // 'd6293
      10'd531  : in_data <= 14'h1867; // 'd6247
      10'd532  : in_data <= 14'h1554; // 'd5460
      10'd533  : in_data <= 14'h0e88; // 'd3720
      10'd534  : in_data <= 14'h07f8; // 'd2040
      10'd535  : in_data <= 14'h121b; // 'd4635
      10'd536  : in_data <= 14'h0a5b; // 'd2651
      10'd537  : in_data <= 14'h080c; // 'd2060
      10'd538  : in_data <= 14'h03b7; // 'd951
      10'd539  : in_data <= 14'h18e4; // 'd6372
      10'd540  : in_data <= 14'h19c1; // 'd6593
      10'd541  : in_data <= 14'h0036; // 'd54
      10'd542  : in_data <= 14'h191d; // 'd6429
      10'd543  : in_data <= 14'h1b14; // 'd6932
      10'd544  : in_data <= 14'h021a; // 'd538
      10'd545  : in_data <= 14'h0528; // 'd1320
      10'd546  : in_data <= 14'h01c3; // 'd451
      10'd547  : in_data <= 14'h0b3c; // 'd2876
      10'd548  : in_data <= 14'h0b4b; // 'd2891
      10'd549  : in_data <= 14'h1673; // 'd5747
      10'd550  : in_data <= 14'h1a5d; // 'd6749
      10'd551  : in_data <= 14'h0237; // 'd567
      10'd552  : in_data <= 14'h036b; // 'd875
      10'd553  : in_data <= 14'h0436; // 'd1078
      10'd554  : in_data <= 14'h1a5a; // 'd6746
      10'd555  : in_data <= 14'h042d; // 'd1069
      10'd556  : in_data <= 14'h0add; // 'd2781
      10'd557  : in_data <= 14'h1090; // 'd4240
      10'd558  : in_data <= 14'h18e6; // 'd6374
      10'd559  : in_data <= 14'h048c; // 'd1164
      10'd560  : in_data <= 14'h1b8b; // 'd7051
      10'd561  : in_data <= 14'h192f; // 'd6447
      10'd562  : in_data <= 14'h1b66; // 'd7014
      10'd563  : in_data <= 14'h0169; // 'd361
      10'd564  : in_data <= 14'h176a; // 'd5994
      10'd565  : in_data <= 14'h0fd7; // 'd4055
      10'd566  : in_data <= 14'h03f2; // 'd1010
      10'd567  : in_data <= 14'h033d; // 'd829
      10'd568  : in_data <= 14'h0351; // 'd849
      10'd569  : in_data <= 14'h15ac; // 'd5548
      10'd570  : in_data <= 14'h01f5; // 'd501
      10'd571  : in_data <= 14'h0d49; // 'd3401
      10'd572  : in_data <= 14'h19aa; // 'd6570
      10'd573  : in_data <= 14'h02ea; // 'd746
      10'd574  : in_data <= 14'h01ef; // 'd495
      10'd575  : in_data <= 14'h05ab; // 'd1451
      10'd576  : in_data <= 14'h078c; // 'd1932
      10'd577  : in_data <= 14'h1153; // 'd4435
      10'd578  : in_data <= 14'h19cb; // 'd6603
      10'd579  : in_data <= 14'h0458; // 'd1112
      10'd580  : in_data <= 14'h107f; // 'd4223
      10'd581  : in_data <= 14'h0b40; // 'd2880
      10'd582  : in_data <= 14'h1152; // 'd4434
      10'd583  : in_data <= 14'h18b2; // 'd6322
      10'd584  : in_data <= 14'h0536; // 'd1334
      10'd585  : in_data <= 14'h1183; // 'd4483
      10'd586  : in_data <= 14'h07bf; // 'd1983
      10'd587  : in_data <= 14'h0e51; // 'd3665
      10'd588  : in_data <= 14'h1652; // 'd5714
      10'd589  : in_data <= 14'h0b98; // 'd2968
      10'd590  : in_data <= 14'h1b92; // 'd7058
      10'd591  : in_data <= 14'h1ba2; // 'd7074
      10'd592  : in_data <= 14'h0462; // 'd1122
      10'd593  : in_data <= 14'h0a8e; // 'd2702
      10'd594  : in_data <= 14'h0b10; // 'd2832
      10'd595  : in_data <= 14'h081a; // 'd2074
      10'd596  : in_data <= 14'h0a6d; // 'd2669
      10'd597  : in_data <= 14'h03d2; // 'd978
      10'd598  : in_data <= 14'h071f; // 'd1823
      10'd599  : in_data <= 14'h0e3b; // 'd3643
      10'd600  : in_data <= 14'h039f; // 'd927
      10'd601  : in_data <= 14'h0dbc; // 'd3516
      10'd602  : in_data <= 14'h1528; // 'd5416
      10'd603  : in_data <= 14'h1219; // 'd4633
      10'd604  : in_data <= 14'h0f1e; // 'd3870
      10'd605  : in_data <= 14'h0828; // 'd2088
      10'd606  : in_data <= 14'h110e; // 'd4366
      10'd607  : in_data <= 14'h12f7; // 'd4855
      10'd608  : in_data <= 14'h16d9; // 'd5849
      10'd609  : in_data <= 14'h1a06; // 'd6662
      10'd610  : in_data <= 14'h0bff; // 'd3071
      10'd611  : in_data <= 14'h0e4a; // 'd3658
      10'd612  : in_data <= 14'h021a; // 'd538
      10'd613  : in_data <= 14'h07de; // 'd2014
      10'd614  : in_data <= 14'h104c; // 'd4172
      10'd615  : in_data <= 14'h0db4; // 'd3508
      10'd616  : in_data <= 14'h11ce; // 'd4558
      10'd617  : in_data <= 14'h0a0d; // 'd2573
      10'd618  : in_data <= 14'h0c66; // 'd3174
      10'd619  : in_data <= 14'h1102; // 'd4354
      10'd620  : in_data <= 14'h10a0; // 'd4256
      10'd621  : in_data <= 14'h18cc; // 'd6348
      10'd622  : in_data <= 14'h1165; // 'd4453
      10'd623  : in_data <= 14'h14f3; // 'd5363
      10'd624  : in_data <= 14'h06a8; // 'd1704
      10'd625  : in_data <= 14'h03c2; // 'd962
      10'd626  : in_data <= 14'h19c6; // 'd6598
      10'd627  : in_data <= 14'h1322; // 'd4898
      10'd628  : in_data <= 14'h10ed; // 'd4333
      10'd629  : in_data <= 14'h0f7c; // 'd3964
      10'd630  : in_data <= 14'h1753; // 'd5971
      10'd631  : in_data <= 14'h0315; // 'd789
      10'd632  : in_data <= 14'h0b30; // 'd2864
      10'd633  : in_data <= 14'h0ff7; // 'd4087
      10'd634  : in_data <= 14'h0d15; // 'd3349
      10'd635  : in_data <= 14'h025f; // 'd607
      10'd636  : in_data <= 14'h1356; // 'd4950
      10'd637  : in_data <= 14'h0a2e; // 'd2606
      10'd638  : in_data <= 14'h0baf; // 'd2991
      10'd639  : in_data <= 14'h12e7; // 'd4839
      10'd640  : in_data <= 14'h01ee; // 'd494
      10'd641  : in_data <= 14'h04fc; // 'd1276
      10'd642  : in_data <= 14'h0322; // 'd802
      10'd643  : in_data <= 14'h16a1; // 'd5793
      10'd644  : in_data <= 14'h05d1; // 'd1489
      10'd645  : in_data <= 14'h1533; // 'd5427
      10'd646  : in_data <= 14'h0f9d; // 'd3997
      10'd647  : in_data <= 14'h129b; // 'd4763
      10'd648  : in_data <= 14'h1216; // 'd4630
      10'd649  : in_data <= 14'h14d5; // 'd5333
      10'd650  : in_data <= 14'h097b; // 'd2427
      10'd651  : in_data <= 14'h0f02; // 'd3842
      10'd652  : in_data <= 14'h0fa0; // 'd4000
      10'd653  : in_data <= 14'h10de; // 'd4318
      10'd654  : in_data <= 14'h1529; // 'd5417
      10'd655  : in_data <= 14'h0487; // 'd1159
      10'd656  : in_data <= 14'h1424; // 'd5156
      10'd657  : in_data <= 14'h1505; // 'd5381
      10'd658  : in_data <= 14'h0192; // 'd402
      10'd659  : in_data <= 14'h1976; // 'd6518
      10'd660  : in_data <= 14'h15ad; // 'd5549
      10'd661  : in_data <= 14'h1ae1; // 'd6881
      10'd662  : in_data <= 14'h108a; // 'd4234
      10'd663  : in_data <= 14'h01ae; // 'd430
      10'd664  : in_data <= 14'h1971; // 'd6513
      10'd665  : in_data <= 14'h16bc; // 'd5820
      10'd666  : in_data <= 14'h08f9; // 'd2297
      10'd667  : in_data <= 14'h0204; // 'd516
      10'd668  : in_data <= 14'h00ad; // 'd173
      10'd669  : in_data <= 14'h014e; // 'd334
      10'd670  : in_data <= 14'h0ec7; // 'd3783
      10'd671  : in_data <= 14'h0a5f; // 'd2655
      10'd672  : in_data <= 14'h19aa; // 'd6570
      10'd673  : in_data <= 14'h0e37; // 'd3639
      10'd674  : in_data <= 14'h1a30; // 'd6704
      10'd675  : in_data <= 14'h0bfe; // 'd3070
      10'd676  : in_data <= 14'h1461; // 'd5217
      10'd677  : in_data <= 14'h13e4; // 'd5092
      10'd678  : in_data <= 14'h1425; // 'd5157
      10'd679  : in_data <= 14'h125a; // 'd4698
      10'd680  : in_data <= 14'h16b1; // 'd5809
      10'd681  : in_data <= 14'h0595; // 'd1429
      10'd682  : in_data <= 14'h12c6; // 'd4806
      10'd683  : in_data <= 14'h0b03; // 'd2819
      10'd684  : in_data <= 14'h1500; // 'd5376
      10'd685  : in_data <= 14'h0b10; // 'd2832
      10'd686  : in_data <= 14'h13fb; // 'd5115
      10'd687  : in_data <= 14'h09c3; // 'd2499
      10'd688  : in_data <= 14'h074e; // 'd1870
      10'd689  : in_data <= 14'h1b11; // 'd6929
      10'd690  : in_data <= 14'h1b8c; // 'd7052
      10'd691  : in_data <= 14'h01d8; // 'd472
      10'd692  : in_data <= 14'h07d7; // 'd2007
      10'd693  : in_data <= 14'h0b65; // 'd2917
      10'd694  : in_data <= 14'h15a2; // 'd5538
      10'd695  : in_data <= 14'h0303; // 'd771
      10'd696  : in_data <= 14'h1b0e; // 'd6926
      10'd697  : in_data <= 14'h1096; // 'd4246
      10'd698  : in_data <= 14'h18e3; // 'd6371
      10'd699  : in_data <= 14'h182a; // 'd6186
      10'd700  : in_data <= 14'h0d31; // 'd3377
      10'd701  : in_data <= 14'h0098; // 'd152
      10'd702  : in_data <= 14'h0a33; // 'd2611
      10'd703  : in_data <= 14'h0b3d; // 'd2877
      10'd704  : in_data <= 14'h05f7; // 'd1527
      10'd705  : in_data <= 14'h07f3; // 'd2035
      10'd706  : in_data <= 14'h08e5; // 'd2277
      10'd707  : in_data <= 14'h044b; // 'd1099
      10'd708  : in_data <= 14'h03e6; // 'd998
      10'd709  : in_data <= 14'h00d0; // 'd208
      10'd710  : in_data <= 14'h0d00; // 'd3328
      10'd711  : in_data <= 14'h0ecf; // 'd3791
      10'd712  : in_data <= 14'h0968; // 'd2408
      10'd713  : in_data <= 14'h0259; // 'd601
      10'd714  : in_data <= 14'h173d; // 'd5949
      10'd715  : in_data <= 14'h1496; // 'd5270
      10'd716  : in_data <= 14'h03c6; // 'd966
      10'd717  : in_data <= 14'h182e; // 'd6190
      10'd718  : in_data <= 14'h17e7; // 'd6119
      10'd719  : in_data <= 14'h0e40; // 'd3648
      10'd720  : in_data <= 14'h0ed1; // 'd3793
      10'd721  : in_data <= 14'h0d96; // 'd3478
      10'd722  : in_data <= 14'h0806; // 'd2054
      10'd723  : in_data <= 14'h0723; // 'd1827
      10'd724  : in_data <= 14'h0736; // 'd1846
      10'd725  : in_data <= 14'h0af2; // 'd2802
      10'd726  : in_data <= 14'h0cfb; // 'd3323
      10'd727  : in_data <= 14'h1092; // 'd4242
      10'd728  : in_data <= 14'h0c90; // 'd3216
      10'd729  : in_data <= 14'h0910; // 'd2320
      10'd730  : in_data <= 14'h05d4; // 'd1492
      10'd731  : in_data <= 14'h05ca; // 'd1482
      10'd732  : in_data <= 14'h0f4c; // 'd3916
      10'd733  : in_data <= 14'h136f; // 'd4975
      10'd734  : in_data <= 14'h0a05; // 'd2565
      10'd735  : in_data <= 14'h17d3; // 'd6099
      10'd736  : in_data <= 14'h1778; // 'd6008
      10'd737  : in_data <= 14'h0859; // 'd2137
      10'd738  : in_data <= 14'h02f3; // 'd755
      10'd739  : in_data <= 14'h14fa; // 'd5370
      10'd740  : in_data <= 14'h0a3b; // 'd2619
      10'd741  : in_data <= 14'h1944; // 'd6468
      10'd742  : in_data <= 14'h0fba; // 'd4026
      10'd743  : in_data <= 14'h0236; // 'd566
      10'd744  : in_data <= 14'h06be; // 'd1726
      10'd745  : in_data <= 14'h04f0; // 'd1264
      10'd746  : in_data <= 14'h1222; // 'd4642
      10'd747  : in_data <= 14'h1b03; // 'd6915
      10'd748  : in_data <= 14'h1780; // 'd6016
      10'd749  : in_data <= 14'h1408; // 'd5128
      10'd750  : in_data <= 14'h041e; // 'd1054
      10'd751  : in_data <= 14'h15cf; // 'd5583
      10'd752  : in_data <= 14'h03aa; // 'd938
      10'd753  : in_data <= 14'h0066; // 'd102
      10'd754  : in_data <= 14'h19ed; // 'd6637
      10'd755  : in_data <= 14'h171b; // 'd5915
      10'd756  : in_data <= 14'h1aae; // 'd6830
      10'd757  : in_data <= 14'h1754; // 'd5972
      10'd758  : in_data <= 14'h0b21; // 'd2849
      10'd759  : in_data <= 14'h0646; // 'd1606
      10'd760  : in_data <= 14'h0055; // 'd85
      10'd761  : in_data <= 14'h04ec; // 'd1260
      10'd762  : in_data <= 14'h0355; // 'd853
      10'd763  : in_data <= 14'h01b7; // 'd439
      10'd764  : in_data <= 14'h052e; // 'd1326
      10'd765  : in_data <= 14'h0070; // 'd112
      10'd766  : in_data <= 14'h0f84; // 'd3972
      10'd767  : in_data <= 14'h0105; // 'd261
      10'd768  : in_data <= 14'h0a9a; // 'd2714
      10'd769  : in_data <= 14'h10a3; // 'd4259
      10'd770  : in_data <= 14'h11ab; // 'd4523
      10'd771  : in_data <= 14'h11fa; // 'd4602
      10'd772  : in_data <= 14'h0045; // 'd69
      10'd773  : in_data <= 14'h19ca; // 'd6602
      10'd774  : in_data <= 14'h187f; // 'd6271
      10'd775  : in_data <= 14'h1371; // 'd4977
      10'd776  : in_data <= 14'h0afc; // 'd2812
      10'd777  : in_data <= 14'h0696; // 'd1686
      10'd778  : in_data <= 14'h1a4a; // 'd6730
      10'd779  : in_data <= 14'h1ab8; // 'd6840
      10'd780  : in_data <= 14'h12de; // 'd4830
      10'd781  : in_data <= 14'h165a; // 'd5722
      10'd782  : in_data <= 14'h03b3; // 'd947
      10'd783  : in_data <= 14'h0aff; // 'd2815
      10'd784  : in_data <= 14'h1a6c; // 'd6764
      10'd785  : in_data <= 14'h048f; // 'd1167
      10'd786  : in_data <= 14'h1752; // 'd5970
      10'd787  : in_data <= 14'h1a1d; // 'd6685
      10'd788  : in_data <= 14'h0ef9; // 'd3833
      10'd789  : in_data <= 14'h0e79; // 'd3705
      10'd790  : in_data <= 14'h18d4; // 'd6356
      10'd791  : in_data <= 14'h07f9; // 'd2041
      10'd792  : in_data <= 14'h1b2a; // 'd6954
      10'd793  : in_data <= 14'h0620; // 'd1568
      10'd794  : in_data <= 14'h0153; // 'd339
      10'd795  : in_data <= 14'h17f2; // 'd6130
      10'd796  : in_data <= 14'h0457; // 'd1111
      10'd797  : in_data <= 14'h16a4; // 'd5796
      10'd798  : in_data <= 14'h055b; // 'd1371
      10'd799  : in_data <= 14'h0bb3; // 'd2995
      10'd800  : in_data <= 14'h18ee; // 'd6382
      10'd801  : in_data <= 14'h1465; // 'd5221
      10'd802  : in_data <= 14'h0cec; // 'd3308
      10'd803  : in_data <= 14'h0775; // 'd1909
      10'd804  : in_data <= 14'h13cd; // 'd5069
      10'd805  : in_data <= 14'h0ec4; // 'd3780
      10'd806  : in_data <= 14'h10ed; // 'd4333
      10'd807  : in_data <= 14'h07a7; // 'd1959
      10'd808  : in_data <= 14'h1174; // 'd4468
      10'd809  : in_data <= 14'h0bc3; // 'd3011
      10'd810  : in_data <= 14'h0aa1; // 'd2721
      10'd811  : in_data <= 14'h16eb; // 'd5867
      10'd812  : in_data <= 14'h0959; // 'd2393
      10'd813  : in_data <= 14'h0f9b; // 'd3995
      10'd814  : in_data <= 14'h1591; // 'd5521
      10'd815  : in_data <= 14'h006e; // 'd110
      10'd816  : in_data <= 14'h1666; // 'd5734
      10'd817  : in_data <= 14'h1b8c; // 'd7052
      10'd818  : in_data <= 14'h1014; // 'd4116
      10'd819  : in_data <= 14'h010d; // 'd269
      10'd820  : in_data <= 14'h135f; // 'd4959
      10'd821  : in_data <= 14'h16f5; // 'd5877
      10'd822  : in_data <= 14'h12ae; // 'd4782
      10'd823  : in_data <= 14'h19ca; // 'd6602
      10'd824  : in_data <= 14'h11d6; // 'd4566
      10'd825  : in_data <= 14'h14bb; // 'd5307
      10'd826  : in_data <= 14'h1a84; // 'd6788
      10'd827  : in_data <= 14'h0d27; // 'd3367
      10'd828  : in_data <= 14'h0f4a; // 'd3914
      10'd829  : in_data <= 14'h08e5; // 'd2277
      10'd830  : in_data <= 14'h056d; // 'd1389
      10'd831  : in_data <= 14'h1708; // 'd5896
      10'd832  : in_data <= 14'h0f3a; // 'd3898
      10'd833  : in_data <= 14'h006b; // 'd107
      10'd834  : in_data <= 14'h1a11; // 'd6673
      10'd835  : in_data <= 14'h0bff; // 'd3071
      10'd836  : in_data <= 14'h1075; // 'd4213
      10'd837  : in_data <= 14'h07b3; // 'd1971
      10'd838  : in_data <= 14'h1326; // 'd4902
      10'd839  : in_data <= 14'h1387; // 'd4999
      10'd840  : in_data <= 14'h0c76; // 'd3190
      10'd841  : in_data <= 14'h139b; // 'd5019
      10'd842  : in_data <= 14'h0abb; // 'd2747
      10'd843  : in_data <= 14'h0e4a; // 'd3658
      10'd844  : in_data <= 14'h19ef; // 'd6639
      10'd845  : in_data <= 14'h07f8; // 'd2040
      10'd846  : in_data <= 14'h00e8; // 'd232
      10'd847  : in_data <= 14'h0b3d; // 'd2877
      10'd848  : in_data <= 14'h126b; // 'd4715
      10'd849  : in_data <= 14'h134c; // 'd4940
      10'd850  : in_data <= 14'h11b7; // 'd4535
      10'd851  : in_data <= 14'h1858; // 'd6232
      10'd852  : in_data <= 14'h0de2; // 'd3554
      10'd853  : in_data <= 14'h173b; // 'd5947
      10'd854  : in_data <= 14'h03c0; // 'd960
      10'd855  : in_data <= 14'h139c; // 'd5020
      10'd856  : in_data <= 14'h0232; // 'd562
      10'd857  : in_data <= 14'h0577; // 'd1399
      10'd858  : in_data <= 14'h1814; // 'd6164
      10'd859  : in_data <= 14'h0c79; // 'd3193
      10'd860  : in_data <= 14'h0c2c; // 'd3116
      10'd861  : in_data <= 14'h1ab7; // 'd6839
      10'd862  : in_data <= 14'h0f78; // 'd3960
      10'd863  : in_data <= 14'h077f; // 'd1919
      10'd864  : in_data <= 14'h129b; // 'd4763
      10'd865  : in_data <= 14'h0b76; // 'd2934
      10'd866  : in_data <= 14'h00ea; // 'd234
      10'd867  : in_data <= 14'h10b2; // 'd4274
      10'd868  : in_data <= 14'h06e2; // 'd1762
      10'd869  : in_data <= 14'h006c; // 'd108
      10'd870  : in_data <= 14'h14e6; // 'd5350
      10'd871  : in_data <= 14'h1416; // 'd5142
      10'd872  : in_data <= 14'h06bc; // 'd1724
      10'd873  : in_data <= 14'h01d5; // 'd469
      10'd874  : in_data <= 14'h152f; // 'd5423
      10'd875  : in_data <= 14'h09be; // 'd2494
      10'd876  : in_data <= 14'h12da; // 'd4826
      10'd877  : in_data <= 14'h0263; // 'd611
      10'd878  : in_data <= 14'h11b3; // 'd4531
      10'd879  : in_data <= 14'h038c; // 'd908
      10'd880  : in_data <= 14'h02f8; // 'd760
      10'd881  : in_data <= 14'h125c; // 'd4700
      10'd882  : in_data <= 14'h188d; // 'd6285
      10'd883  : in_data <= 14'h054e; // 'd1358
      10'd884  : in_data <= 14'h1509; // 'd5385
      10'd885  : in_data <= 14'h19f7; // 'd6647
      10'd886  : in_data <= 14'h0906; // 'd2310
      10'd887  : in_data <= 14'h0eac; // 'd3756
      10'd888  : in_data <= 14'h1106; // 'd4358
      10'd889  : in_data <= 14'h1296; // 'd4758
      10'd890  : in_data <= 14'h0e24; // 'd3620
      10'd891  : in_data <= 14'h10fe; // 'd4350
      10'd892  : in_data <= 14'h17f1; // 'd6129
      10'd893  : in_data <= 14'h13a5; // 'd5029
      10'd894  : in_data <= 14'h1186; // 'd4486
      10'd895  : in_data <= 14'h1229; // 'd4649
      10'd896  : in_data <= 14'h05d5; // 'd1493
      10'd897  : in_data <= 14'h00ce; // 'd206
      10'd898  : in_data <= 14'h0f53; // 'd3923
      10'd899  : in_data <= 14'h02fd; // 'd765
      10'd900  : in_data <= 14'h1b33; // 'd6963
      10'd901  : in_data <= 14'h1010; // 'd4112
      10'd902  : in_data <= 14'h1a1d; // 'd6685
      10'd903  : in_data <= 14'h172f; // 'd5935
      10'd904  : in_data <= 14'h12ae; // 'd4782
      10'd905  : in_data <= 14'h0fb0; // 'd4016
      10'd906  : in_data <= 14'h0639; // 'd1593
      10'd907  : in_data <= 14'h08c2; // 'd2242
      10'd908  : in_data <= 14'h177e; // 'd6014
      10'd909  : in_data <= 14'h0495; // 'd1173
      10'd910  : in_data <= 14'h1473; // 'd5235
      10'd911  : in_data <= 14'h0e60; // 'd3680
      10'd912  : in_data <= 14'h0479; // 'd1145
      10'd913  : in_data <= 14'h0a0f; // 'd2575
      10'd914  : in_data <= 14'h08b6; // 'd2230
      10'd915  : in_data <= 14'h0d1c; // 'd3356
      10'd916  : in_data <= 14'h0636; // 'd1590
      10'd917  : in_data <= 14'h07ff; // 'd2047
      10'd918  : in_data <= 14'h10f4; // 'd4340
      10'd919  : in_data <= 14'h0af7; // 'd2807
      10'd920  : in_data <= 14'h1125; // 'd4389
      10'd921  : in_data <= 14'h0a9e; // 'd2718
      10'd922  : in_data <= 14'h1551; // 'd5457
      10'd923  : in_data <= 14'h1508; // 'd5384
      10'd924  : in_data <= 14'h0b37; // 'd2871
      10'd925  : in_data <= 14'h139a; // 'd5018
      10'd926  : in_data <= 14'h12d4; // 'd4820
      10'd927  : in_data <= 14'h19ff; // 'd6655
      10'd928  : in_data <= 14'h1409; // 'd5129
      10'd929  : in_data <= 14'h1526; // 'd5414
      10'd930  : in_data <= 14'h0658; // 'd1624
      10'd931  : in_data <= 14'h11c7; // 'd4551
      10'd932  : in_data <= 14'h1094; // 'd4244
      10'd933  : in_data <= 14'h10d8; // 'd4312
      10'd934  : in_data <= 14'h0c62; // 'd3170
      10'd935  : in_data <= 14'h032b; // 'd811
      10'd936  : in_data <= 14'h1601; // 'd5633
      10'd937  : in_data <= 14'h060d; // 'd1549
      10'd938  : in_data <= 14'h179c; // 'd6044
      10'd939  : in_data <= 14'h14a2; // 'd5282
      10'd940  : in_data <= 14'h0479; // 'd1145
      10'd941  : in_data <= 14'h0a26; // 'd2598
      10'd942  : in_data <= 14'h0ce2; // 'd3298
      10'd943  : in_data <= 14'h1989; // 'd6537
      10'd944  : in_data <= 14'h1af1; // 'd6897
      10'd945  : in_data <= 14'h0637; // 'd1591
      10'd946  : in_data <= 14'h058b; // 'd1419
      10'd947  : in_data <= 14'h0030; // 'd48
      10'd948  : in_data <= 14'h0429; // 'd1065
      10'd949  : in_data <= 14'h02ed; // 'd749
      10'd950  : in_data <= 14'h0ef4; // 'd3828
      10'd951  : in_data <= 14'h0a3b; // 'd2619
      10'd952  : in_data <= 14'h1879; // 'd6265
      10'd953  : in_data <= 14'h16fa; // 'd5882
      10'd954  : in_data <= 14'h08ff; // 'd2303
      10'd955  : in_data <= 14'h0a97; // 'd2711
      10'd956  : in_data <= 14'h1128; // 'd4392
      10'd957  : in_data <= 14'h113b; // 'd4411
      10'd958  : in_data <= 14'h12a4; // 'd4772
      10'd959  : in_data <= 14'h16ec; // 'd5868
      10'd960  : in_data <= 14'h0c10; // 'd3088
      10'd961  : in_data <= 14'h0c72; // 'd3186
      10'd962  : in_data <= 14'h0939; // 'd2361
      10'd963  : in_data <= 14'h109c; // 'd4252
      10'd964  : in_data <= 14'h0beb; // 'd3051
      10'd965  : in_data <= 14'h0476; // 'd1142
      10'd966  : in_data <= 14'h0772; // 'd1906
      10'd967  : in_data <= 14'h1215; // 'd4629
      10'd968  : in_data <= 14'h1421; // 'd5153
      10'd969  : in_data <= 14'h06a5; // 'd1701
      10'd970  : in_data <= 14'h0900; // 'd2304
      10'd971  : in_data <= 14'h17a5; // 'd6053
      10'd972  : in_data <= 14'h1520; // 'd5408
      10'd973  : in_data <= 14'h032b; // 'd811
      10'd974  : in_data <= 14'h0ce2; // 'd3298
      10'd975  : in_data <= 14'h10ca; // 'd4298
      10'd976  : in_data <= 14'h0c1f; // 'd3103
      10'd977  : in_data <= 14'h015f; // 'd351
      10'd978  : in_data <= 14'h0770; // 'd1904
      10'd979  : in_data <= 14'h1aba; // 'd6842
      10'd980  : in_data <= 14'h1946; // 'd6470
      10'd981  : in_data <= 14'h1762; // 'd5986
      10'd982  : in_data <= 14'h092b; // 'd2347
      10'd983  : in_data <= 14'h0e30; // 'd3632
      10'd984  : in_data <= 14'h1999; // 'd6553
      10'd985  : in_data <= 14'h157c; // 'd5500
      10'd986  : in_data <= 14'h095e; // 'd2398
      10'd987  : in_data <= 14'h02a8; // 'd680
      10'd988  : in_data <= 14'h04e2; // 'd1250
      10'd989  : in_data <= 14'h002d; // 'd45
      10'd990  : in_data <= 14'h0adc; // 'd2780
      10'd991  : in_data <= 14'h1157; // 'd4439
      10'd992  : in_data <= 14'h145c; // 'd5212
      10'd993  : in_data <= 14'h1446; // 'd5190
      10'd994  : in_data <= 14'h1520; // 'd5408
      10'd995  : in_data <= 14'h028c; // 'd652
      10'd996  : in_data <= 14'h04fc; // 'd1276
      10'd997  : in_data <= 14'h14c7; // 'd5319
      10'd998  : in_data <= 14'h0e19; // 'd3609
      10'd999  : in_data <= 14'h06bc; // 'd1724
      10'd1000 : in_data <= 14'h1c02; // 'd7170
      10'd1001 : in_data <= 14'h199e; // 'd6558
      10'd1002 : in_data <= 14'h1983; // 'd6531
      10'd1003 : in_data <= 14'h1178; // 'd4472
      10'd1004 : in_data <= 14'h1627; // 'd5671
      10'd1005 : in_data <= 14'h11f4; // 'd4596
      10'd1006 : in_data <= 14'h067a; // 'd1658
      10'd1007 : in_data <= 14'h0ca0; // 'd3232
      10'd1008 : in_data <= 14'h155b; // 'd5467
      10'd1009 : in_data <= 14'h1528; // 'd5416
      10'd1010 : in_data <= 14'h0245; // 'd581
      10'd1011 : in_data <= 14'h03b5; // 'd949
      10'd1012 : in_data <= 14'h0788; // 'd1928
      default  : in_data <= 14'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      11'd0    : out_data_ref <= 8'h30;
      11'd1    : out_data_ref <= 8'h46;
      11'd2    : out_data_ref <= 8'hec;
      11'd3    : out_data_ref <= 8'h85;
      11'd4    : out_data_ref <= 8'hb9;
      11'd5    : out_data_ref <= 8'hde;
      11'd6    : out_data_ref <= 8'h48;
      11'd7    : out_data_ref <= 8'h1f;
      11'd8    : out_data_ref <= 8'hae;
      11'd9    : out_data_ref <= 8'hbf;
      11'd10   : out_data_ref <= 8'h95;
      11'd11   : out_data_ref <= 8'hd1;
      11'd12   : out_data_ref <= 8'h9b;
      11'd13   : out_data_ref <= 8'hba;
      11'd14   : out_data_ref <= 8'h38;
      11'd15   : out_data_ref <= 8'hfd;
      11'd16   : out_data_ref <= 8'heb;
      11'd17   : out_data_ref <= 8'ha9;
      11'd18   : out_data_ref <= 8'he8;
      11'd19   : out_data_ref <= 8'heb;
      11'd20   : out_data_ref <= 8'hed;
      11'd21   : out_data_ref <= 8'h54;
      11'd22   : out_data_ref <= 8'hdd;
      11'd23   : out_data_ref <= 8'h01;
      11'd24   : out_data_ref <= 8'haa;
      11'd25   : out_data_ref <= 8'h79;
      11'd26   : out_data_ref <= 8'h54;
      11'd27   : out_data_ref <= 8'h04;
      11'd28   : out_data_ref <= 8'hba;
      11'd29   : out_data_ref <= 8'h11;
      11'd30   : out_data_ref <= 8'h27;
      11'd31   : out_data_ref <= 8'h60;
      11'd32   : out_data_ref <= 8'h94;
      11'd33   : out_data_ref <= 8'hd1;
      11'd34   : out_data_ref <= 8'hf6;
      11'd35   : out_data_ref <= 8'hf9;
      11'd36   : out_data_ref <= 8'h99;
      11'd37   : out_data_ref <= 8'hff;
      11'd38   : out_data_ref <= 8'h9e;
      11'd39   : out_data_ref <= 8'h27;
      11'd40   : out_data_ref <= 8'h92;
      11'd41   : out_data_ref <= 8'h00;
      11'd42   : out_data_ref <= 8'hb0;
      11'd43   : out_data_ref <= 8'h67;
      11'd44   : out_data_ref <= 8'hb6;
      11'd45   : out_data_ref <= 8'h4c;
      11'd46   : out_data_ref <= 8'h17;
      11'd47   : out_data_ref <= 8'hea;
      11'd48   : out_data_ref <= 8'hc8;
      11'd49   : out_data_ref <= 8'ha6;
      11'd50   : out_data_ref <= 8'h30;
      11'd51   : out_data_ref <= 8'h33;
      11'd52   : out_data_ref <= 8'hdc;
      11'd53   : out_data_ref <= 8'h6e;
      11'd54   : out_data_ref <= 8'hd5;
      11'd55   : out_data_ref <= 8'h75;
      11'd56   : out_data_ref <= 8'hb1;
      11'd57   : out_data_ref <= 8'h20;
      11'd58   : out_data_ref <= 8'h45;
      11'd59   : out_data_ref <= 8'h0a;
      11'd60   : out_data_ref <= 8'hdc;
      11'd61   : out_data_ref <= 8'ha5;
      11'd62   : out_data_ref <= 8'h45;
      11'd63   : out_data_ref <= 8'h06;
      11'd64   : out_data_ref <= 8'h74;
      11'd65   : out_data_ref <= 8'h55;
      11'd66   : out_data_ref <= 8'h41;
      11'd67   : out_data_ref <= 8'h50;
      11'd68   : out_data_ref <= 8'h9e;
      11'd69   : out_data_ref <= 8'h4e;
      11'd70   : out_data_ref <= 8'h18;
      11'd71   : out_data_ref <= 8'h24;
      11'd72   : out_data_ref <= 8'hd5;
      11'd73   : out_data_ref <= 8'h22;
      11'd74   : out_data_ref <= 8'hfb;
      11'd75   : out_data_ref <= 8'hfc;
      11'd76   : out_data_ref <= 8'h3f;
      11'd77   : out_data_ref <= 8'hb2;
      11'd78   : out_data_ref <= 8'h9e;
      11'd79   : out_data_ref <= 8'hc7;
      11'd80   : out_data_ref <= 8'h86;
      11'd81   : out_data_ref <= 8'ha1;
      11'd82   : out_data_ref <= 8'h90;
      11'd83   : out_data_ref <= 8'h12;
      11'd84   : out_data_ref <= 8'haa;
      11'd85   : out_data_ref <= 8'h80;
      11'd86   : out_data_ref <= 8'h15;
      11'd87   : out_data_ref <= 8'h16;
      11'd88   : out_data_ref <= 8'h44;
      11'd89   : out_data_ref <= 8'h6b;
      11'd90   : out_data_ref <= 8'h06;
      11'd91   : out_data_ref <= 8'he0;
      11'd92   : out_data_ref <= 8'hdd;
      11'd93   : out_data_ref <= 8'h23;
      11'd94   : out_data_ref <= 8'h9b;
      11'd95   : out_data_ref <= 8'he6;
      11'd96   : out_data_ref <= 8'hd4;
      11'd97   : out_data_ref <= 8'h6d;
      11'd98   : out_data_ref <= 8'h13;
      11'd99   : out_data_ref <= 8'hc0;
      11'd100  : out_data_ref <= 8'hc3;
      11'd101  : out_data_ref <= 8'hff;
      11'd102  : out_data_ref <= 8'h30;
      11'd103  : out_data_ref <= 8'h30;
      11'd104  : out_data_ref <= 8'h23;
      11'd105  : out_data_ref <= 8'h25;
      11'd106  : out_data_ref <= 8'hf6;
      11'd107  : out_data_ref <= 8'he0;
      11'd108  : out_data_ref <= 8'he1;
      11'd109  : out_data_ref <= 8'h10;
      11'd110  : out_data_ref <= 8'haa;
      11'd111  : out_data_ref <= 8'h71;
      11'd112  : out_data_ref <= 8'hcb;
      11'd113  : out_data_ref <= 8'h49;
      11'd114  : out_data_ref <= 8'h53;
      11'd115  : out_data_ref <= 8'h0b;
      11'd116  : out_data_ref <= 8'h50;
      11'd117  : out_data_ref <= 8'h27;
      11'd118  : out_data_ref <= 8'he1;
      11'd119  : out_data_ref <= 8'h95;
      11'd120  : out_data_ref <= 8'h48;
      11'd121  : out_data_ref <= 8'heb;
      11'd122  : out_data_ref <= 8'hf1;
      11'd123  : out_data_ref <= 8'hb2;
      11'd124  : out_data_ref <= 8'ha6;
      11'd125  : out_data_ref <= 8'h64;
      11'd126  : out_data_ref <= 8'hd6;
      11'd127  : out_data_ref <= 8'hbf;
      11'd128  : out_data_ref <= 8'hc7;
      11'd129  : out_data_ref <= 8'h7e;
      11'd130  : out_data_ref <= 8'h7c;
      11'd131  : out_data_ref <= 8'h3b;
      11'd132  : out_data_ref <= 8'hed;
      11'd133  : out_data_ref <= 8'h1c;
      11'd134  : out_data_ref <= 8'h18;
      11'd135  : out_data_ref <= 8'he0;
      11'd136  : out_data_ref <= 8'he8;
      11'd137  : out_data_ref <= 8'h27;
      11'd138  : out_data_ref <= 8'h08;
      11'd139  : out_data_ref <= 8'h84;
      11'd140  : out_data_ref <= 8'he2;
      11'd141  : out_data_ref <= 8'hdf;
      11'd142  : out_data_ref <= 8'h85;
      11'd143  : out_data_ref <= 8'h3b;
      11'd144  : out_data_ref <= 8'h41;
      11'd145  : out_data_ref <= 8'h6f;
      11'd146  : out_data_ref <= 8'h03;
      11'd147  : out_data_ref <= 8'h60;
      11'd148  : out_data_ref <= 8'h6d;
      11'd149  : out_data_ref <= 8'h1e;
      11'd150  : out_data_ref <= 8'h02;
      11'd151  : out_data_ref <= 8'h93;
      11'd152  : out_data_ref <= 8'he5;
      11'd153  : out_data_ref <= 8'h99;
      11'd154  : out_data_ref <= 8'hb8;
      11'd155  : out_data_ref <= 8'hac;
      11'd156  : out_data_ref <= 8'hc4;
      11'd157  : out_data_ref <= 8'h36;
      11'd158  : out_data_ref <= 8'h40;
      11'd159  : out_data_ref <= 8'h65;
      11'd160  : out_data_ref <= 8'hc5;
      11'd161  : out_data_ref <= 8'h3f;
      11'd162  : out_data_ref <= 8'hed;
      11'd163  : out_data_ref <= 8'hbf;
      11'd164  : out_data_ref <= 8'h1f;
      11'd165  : out_data_ref <= 8'h4f;
      11'd166  : out_data_ref <= 8'h39;
      11'd167  : out_data_ref <= 8'haa;
      11'd168  : out_data_ref <= 8'h70;
      11'd169  : out_data_ref <= 8'h9b;
      11'd170  : out_data_ref <= 8'h7b;
      11'd171  : out_data_ref <= 8'h55;
      11'd172  : out_data_ref <= 8'h31;
      11'd173  : out_data_ref <= 8'hcb;
      11'd174  : out_data_ref <= 8'hf7;
      11'd175  : out_data_ref <= 8'h98;
      11'd176  : out_data_ref <= 8'h0f;
      11'd177  : out_data_ref <= 8'h6e;
      11'd178  : out_data_ref <= 8'h48;
      11'd179  : out_data_ref <= 8'he6;
      11'd180  : out_data_ref <= 8'hd3;
      11'd181  : out_data_ref <= 8'h59;
      11'd182  : out_data_ref <= 8'h4e;
      11'd183  : out_data_ref <= 8'h58;
      11'd184  : out_data_ref <= 8'h87;
      11'd185  : out_data_ref <= 8'h20;
      11'd186  : out_data_ref <= 8'h58;
      11'd187  : out_data_ref <= 8'hdd;
      11'd188  : out_data_ref <= 8'h58;
      11'd189  : out_data_ref <= 8'hb8;
      11'd190  : out_data_ref <= 8'h0c;
      11'd191  : out_data_ref <= 8'h9f;
      11'd192  : out_data_ref <= 8'h3c;
      11'd193  : out_data_ref <= 8'h8c;
      11'd194  : out_data_ref <= 8'h3e;
      11'd195  : out_data_ref <= 8'ha0;
      11'd196  : out_data_ref <= 8'h5f;
      11'd197  : out_data_ref <= 8'h08;
      11'd198  : out_data_ref <= 8'h74;
      11'd199  : out_data_ref <= 8'hec;
      11'd200  : out_data_ref <= 8'h81;
      11'd201  : out_data_ref <= 8'h77;
      11'd202  : out_data_ref <= 8'h4f;
      11'd203  : out_data_ref <= 8'h62;
      11'd204  : out_data_ref <= 8'h29;
      11'd205  : out_data_ref <= 8'h2c;
      11'd206  : out_data_ref <= 8'h12;
      11'd207  : out_data_ref <= 8'h2f;
      11'd208  : out_data_ref <= 8'h13;
      11'd209  : out_data_ref <= 8'h86;
      11'd210  : out_data_ref <= 8'hbd;
      11'd211  : out_data_ref <= 8'hae;
      11'd212  : out_data_ref <= 8'h52;
      11'd213  : out_data_ref <= 8'h19;
      11'd214  : out_data_ref <= 8'ha7;
      11'd215  : out_data_ref <= 8'h64;
      11'd216  : out_data_ref <= 8'h4f;
      11'd217  : out_data_ref <= 8'h39;
      11'd218  : out_data_ref <= 8'hdc;
      11'd219  : out_data_ref <= 8'h56;
      11'd220  : out_data_ref <= 8'h17;
      11'd221  : out_data_ref <= 8'hba;
      11'd222  : out_data_ref <= 8'hfd;
      11'd223  : out_data_ref <= 8'h35;
      11'd224  : out_data_ref <= 8'h2a;
      11'd225  : out_data_ref <= 8'h32;
      11'd226  : out_data_ref <= 8'ha3;
      11'd227  : out_data_ref <= 8'he7;
      11'd228  : out_data_ref <= 8'hd4;
      11'd229  : out_data_ref <= 8'h9f;
      11'd230  : out_data_ref <= 8'h2b;
      11'd231  : out_data_ref <= 8'hcd;
      11'd232  : out_data_ref <= 8'hf9;
      11'd233  : out_data_ref <= 8'hb0;
      11'd234  : out_data_ref <= 8'h68;
      11'd235  : out_data_ref <= 8'hc1;
      11'd236  : out_data_ref <= 8'h3d;
      11'd237  : out_data_ref <= 8'hf7;
      11'd238  : out_data_ref <= 8'h71;
      11'd239  : out_data_ref <= 8'he2;
      11'd240  : out_data_ref <= 8'h84;
      11'd241  : out_data_ref <= 8'h4b;
      11'd242  : out_data_ref <= 8'h56;
      11'd243  : out_data_ref <= 8'he7;
      11'd244  : out_data_ref <= 8'h15;
      11'd245  : out_data_ref <= 8'h1b;
      11'd246  : out_data_ref <= 8'hb3;
      11'd247  : out_data_ref <= 8'h08;
      11'd248  : out_data_ref <= 8'h09;
      11'd249  : out_data_ref <= 8'h37;
      11'd250  : out_data_ref <= 8'hd5;
      11'd251  : out_data_ref <= 8'haf;
      11'd252  : out_data_ref <= 8'h49;
      11'd253  : out_data_ref <= 8'h7e;
      11'd254  : out_data_ref <= 8'h06;
      11'd255  : out_data_ref <= 8'h42;
      11'd256  : out_data_ref <= 8'h64;
      11'd257  : out_data_ref <= 8'hc8;
      11'd258  : out_data_ref <= 8'ha0;
      11'd259  : out_data_ref <= 8'h67;
      11'd260  : out_data_ref <= 8'h94;
      11'd261  : out_data_ref <= 8'h68;
      11'd262  : out_data_ref <= 8'h97;
      11'd263  : out_data_ref <= 8'ha9;
      11'd264  : out_data_ref <= 8'h9c;
      11'd265  : out_data_ref <= 8'h0a;
      11'd266  : out_data_ref <= 8'hfd;
      11'd267  : out_data_ref <= 8'hf3;
      11'd268  : out_data_ref <= 8'h21;
      11'd269  : out_data_ref <= 8'h77;
      11'd270  : out_data_ref <= 8'hc5;
      11'd271  : out_data_ref <= 8'h8c;
      11'd272  : out_data_ref <= 8'h90;
      11'd273  : out_data_ref <= 8'h84;
      11'd274  : out_data_ref <= 8'h9d;
      11'd275  : out_data_ref <= 8'h2f;
      11'd276  : out_data_ref <= 8'hc2;
      11'd277  : out_data_ref <= 8'h7c;
      11'd278  : out_data_ref <= 8'hc7;
      11'd279  : out_data_ref <= 8'hef;
      11'd280  : out_data_ref <= 8'h1f;
      11'd281  : out_data_ref <= 8'h38;
      11'd282  : out_data_ref <= 8'h05;
      11'd283  : out_data_ref <= 8'h62;
      11'd284  : out_data_ref <= 8'h6a;
      11'd285  : out_data_ref <= 8'h58;
      11'd286  : out_data_ref <= 8'h8f;
      11'd287  : out_data_ref <= 8'hb7;
      11'd288  : out_data_ref <= 8'h14;
      11'd289  : out_data_ref <= 8'h67;
      11'd290  : out_data_ref <= 8'h2f;
      11'd291  : out_data_ref <= 8'h8e;
      11'd292  : out_data_ref <= 8'h7e;
      11'd293  : out_data_ref <= 8'h54;
      11'd294  : out_data_ref <= 8'he0;
      11'd295  : out_data_ref <= 8'h5f;
      11'd296  : out_data_ref <= 8'he0;
      11'd297  : out_data_ref <= 8'h11;
      11'd298  : out_data_ref <= 8'hfe;
      11'd299  : out_data_ref <= 8'h69;
      11'd300  : out_data_ref <= 8'h18;
      11'd301  : out_data_ref <= 8'hbd;
      11'd302  : out_data_ref <= 8'hab;
      11'd303  : out_data_ref <= 8'h7e;
      11'd304  : out_data_ref <= 8'he2;
      11'd305  : out_data_ref <= 8'hac;
      11'd306  : out_data_ref <= 8'hb1;
      11'd307  : out_data_ref <= 8'hd6;
      11'd308  : out_data_ref <= 8'h58;
      11'd309  : out_data_ref <= 8'hb8;
      11'd310  : out_data_ref <= 8'hcb;
      11'd311  : out_data_ref <= 8'h9a;
      11'd312  : out_data_ref <= 8'h9a;
      11'd313  : out_data_ref <= 8'hb6;
      11'd314  : out_data_ref <= 8'h46;
      11'd315  : out_data_ref <= 8'hec;
      11'd316  : out_data_ref <= 8'he3;
      11'd317  : out_data_ref <= 8'h45;
      11'd318  : out_data_ref <= 8'h61;
      11'd319  : out_data_ref <= 8'hb1;
      11'd320  : out_data_ref <= 8'h36;
      11'd321  : out_data_ref <= 8'hbb;
      11'd322  : out_data_ref <= 8'hee;
      11'd323  : out_data_ref <= 8'h43;
      11'd324  : out_data_ref <= 8'h61;
      11'd325  : out_data_ref <= 8'hbb;
      11'd326  : out_data_ref <= 8'hfb;
      11'd327  : out_data_ref <= 8'h57;
      11'd328  : out_data_ref <= 8'hce;
      11'd329  : out_data_ref <= 8'h62;
      11'd330  : out_data_ref <= 8'ha4;
      11'd331  : out_data_ref <= 8'h59;
      11'd332  : out_data_ref <= 8'h43;
      11'd333  : out_data_ref <= 8'hf3;
      11'd334  : out_data_ref <= 8'h98;
      11'd335  : out_data_ref <= 8'h43;
      11'd336  : out_data_ref <= 8'h49;
      11'd337  : out_data_ref <= 8'h76;
      11'd338  : out_data_ref <= 8'h13;
      11'd339  : out_data_ref <= 8'h19;
      11'd340  : out_data_ref <= 8'he9;
      11'd341  : out_data_ref <= 8'h01;
      11'd342  : out_data_ref <= 8'hd5;
      11'd343  : out_data_ref <= 8'hfe;
      11'd344  : out_data_ref <= 8'hf3;
      11'd345  : out_data_ref <= 8'hda;
      11'd346  : out_data_ref <= 8'hf0;
      11'd347  : out_data_ref <= 8'hbd;
      11'd348  : out_data_ref <= 8'hb8;
      11'd349  : out_data_ref <= 8'h2d;
      11'd350  : out_data_ref <= 8'h0b;
      11'd351  : out_data_ref <= 8'hdc;
      11'd352  : out_data_ref <= 8'hbd;
      11'd353  : out_data_ref <= 8'h2b;
      11'd354  : out_data_ref <= 8'hc0;
      11'd355  : out_data_ref <= 8'h11;
      11'd356  : out_data_ref <= 8'h54;
      11'd357  : out_data_ref <= 8'hf4;
      11'd358  : out_data_ref <= 8'hf1;
      11'd359  : out_data_ref <= 8'h43;
      11'd360  : out_data_ref <= 8'ha8;
      11'd361  : out_data_ref <= 8'h06;
      11'd362  : out_data_ref <= 8'h3a;
      11'd363  : out_data_ref <= 8'h2c;
      11'd364  : out_data_ref <= 8'hbe;
      11'd365  : out_data_ref <= 8'hd9;
      11'd366  : out_data_ref <= 8'hc2;
      11'd367  : out_data_ref <= 8'hf9;
      11'd368  : out_data_ref <= 8'hed;
      11'd369  : out_data_ref <= 8'h9c;
      11'd370  : out_data_ref <= 8'hc0;
      11'd371  : out_data_ref <= 8'h61;
      11'd372  : out_data_ref <= 8'h85;
      11'd373  : out_data_ref <= 8'h20;
      11'd374  : out_data_ref <= 8'h7f;
      11'd375  : out_data_ref <= 8'h15;
      11'd376  : out_data_ref <= 8'ha3;
      11'd377  : out_data_ref <= 8'h12;
      11'd378  : out_data_ref <= 8'h89;
      11'd379  : out_data_ref <= 8'hf0;
      11'd380  : out_data_ref <= 8'h73;
      11'd381  : out_data_ref <= 8'h56;
      11'd382  : out_data_ref <= 8'h20;
      11'd383  : out_data_ref <= 8'hd2;
      11'd384  : out_data_ref <= 8'hd7;
      11'd385  : out_data_ref <= 8'h1d;
      11'd386  : out_data_ref <= 8'h3e;
      11'd387  : out_data_ref <= 8'hec;
      11'd388  : out_data_ref <= 8'h56;
      11'd389  : out_data_ref <= 8'h16;
      11'd390  : out_data_ref <= 8'h87;
      11'd391  : out_data_ref <= 8'h21;
      11'd392  : out_data_ref <= 8'h0d;
      11'd393  : out_data_ref <= 8'h6a;
      11'd394  : out_data_ref <= 8'h52;
      11'd395  : out_data_ref <= 8'h95;
      11'd396  : out_data_ref <= 8'hdd;
      11'd397  : out_data_ref <= 8'hd9;
      11'd398  : out_data_ref <= 8'h1d;
      11'd399  : out_data_ref <= 8'h46;
      11'd400  : out_data_ref <= 8'h5f;
      11'd401  : out_data_ref <= 8'h8e;
      11'd402  : out_data_ref <= 8'h34;
      11'd403  : out_data_ref <= 8'hd2;
      11'd404  : out_data_ref <= 8'hdd;
      11'd405  : out_data_ref <= 8'h21;
      11'd406  : out_data_ref <= 8'hc4;
      11'd407  : out_data_ref <= 8'h03;
      11'd408  : out_data_ref <= 8'ha5;
      11'd409  : out_data_ref <= 8'h2e;
      11'd410  : out_data_ref <= 8'hc3;
      11'd411  : out_data_ref <= 8'h01;
      11'd412  : out_data_ref <= 8'h33;
      11'd413  : out_data_ref <= 8'h9c;
      11'd414  : out_data_ref <= 8'h1e;
      11'd415  : out_data_ref <= 8'h81;
      11'd416  : out_data_ref <= 8'h11;
      11'd417  : out_data_ref <= 8'hac;
      11'd418  : out_data_ref <= 8'hac;
      11'd419  : out_data_ref <= 8'he4;
      11'd420  : out_data_ref <= 8'h35;
      11'd421  : out_data_ref <= 8'h01;
      11'd422  : out_data_ref <= 8'h33;
      11'd423  : out_data_ref <= 8'h47;
      11'd424  : out_data_ref <= 8'hb4;
      11'd425  : out_data_ref <= 8'h29;
      11'd426  : out_data_ref <= 8'h39;
      11'd427  : out_data_ref <= 8'h8e;
      11'd428  : out_data_ref <= 8'h7f;
      11'd429  : out_data_ref <= 8'hd7;
      11'd430  : out_data_ref <= 8'h0b;
      11'd431  : out_data_ref <= 8'h35;
      11'd432  : out_data_ref <= 8'h74;
      11'd433  : out_data_ref <= 8'h00;
      11'd434  : out_data_ref <= 8'h96;
      11'd435  : out_data_ref <= 8'hdf;
      11'd436  : out_data_ref <= 8'h62;
      11'd437  : out_data_ref <= 8'hb8;
      11'd438  : out_data_ref <= 8'hbd;
      11'd439  : out_data_ref <= 8'h17;
      11'd440  : out_data_ref <= 8'hbf;
      11'd441  : out_data_ref <= 8'hf0;
      11'd442  : out_data_ref <= 8'hc0;
      11'd443  : out_data_ref <= 8'h3b;
      11'd444  : out_data_ref <= 8'ha2;
      11'd445  : out_data_ref <= 8'hf0;
      11'd446  : out_data_ref <= 8'h1e;
      11'd447  : out_data_ref <= 8'hc9;
      11'd448  : out_data_ref <= 8'h27;
      11'd449  : out_data_ref <= 8'h1e;
      11'd450  : out_data_ref <= 8'h25;
      11'd451  : out_data_ref <= 8'h06;
      11'd452  : out_data_ref <= 8'hcf;
      11'd453  : out_data_ref <= 8'h57;
      11'd454  : out_data_ref <= 8'h4f;
      11'd455  : out_data_ref <= 8'h3a;
      11'd456  : out_data_ref <= 8'hc1;
      11'd457  : out_data_ref <= 8'hb3;
      11'd458  : out_data_ref <= 8'h9b;
      11'd459  : out_data_ref <= 8'h23;
      11'd460  : out_data_ref <= 8'h69;
      11'd461  : out_data_ref <= 8'h63;
      11'd462  : out_data_ref <= 8'he8;
      11'd463  : out_data_ref <= 8'h85;
      11'd464  : out_data_ref <= 8'hbc;
      11'd465  : out_data_ref <= 8'h35;
      11'd466  : out_data_ref <= 8'hae;
      11'd467  : out_data_ref <= 8'h7e;
      11'd468  : out_data_ref <= 8'he2;
      11'd469  : out_data_ref <= 8'h85;
      11'd470  : out_data_ref <= 8'hf0;
      11'd471  : out_data_ref <= 8'hea;
      11'd472  : out_data_ref <= 8'h28;
      11'd473  : out_data_ref <= 8'hfe;
      11'd474  : out_data_ref <= 8'hac;
      11'd475  : out_data_ref <= 8'hd7;
      11'd476  : out_data_ref <= 8'h79;
      11'd477  : out_data_ref <= 8'hab;
      11'd478  : out_data_ref <= 8'h22;
      11'd479  : out_data_ref <= 8'h46;
      11'd480  : out_data_ref <= 8'h5f;
      11'd481  : out_data_ref <= 8'h78;
      11'd482  : out_data_ref <= 8'h08;
      11'd483  : out_data_ref <= 8'h9c;
      11'd484  : out_data_ref <= 8'h77;
      11'd485  : out_data_ref <= 8'hc1;
      11'd486  : out_data_ref <= 8'heb;
      11'd487  : out_data_ref <= 8'ha9;
      11'd488  : out_data_ref <= 8'hb2;
      11'd489  : out_data_ref <= 8'h5a;
      11'd490  : out_data_ref <= 8'h85;
      11'd491  : out_data_ref <= 8'hde;
      11'd492  : out_data_ref <= 8'he5;
      11'd493  : out_data_ref <= 8'hf6;
      11'd494  : out_data_ref <= 8'hd7;
      11'd495  : out_data_ref <= 8'h61;
      11'd496  : out_data_ref <= 8'he1;
      11'd497  : out_data_ref <= 8'hc1;
      11'd498  : out_data_ref <= 8'h97;
      11'd499  : out_data_ref <= 8'haf;
      11'd500  : out_data_ref <= 8'h29;
      11'd501  : out_data_ref <= 8'h89;
      11'd502  : out_data_ref <= 8'h81;
      11'd503  : out_data_ref <= 8'hb6;
      11'd504  : out_data_ref <= 8'h88;
      11'd505  : out_data_ref <= 8'h49;
      11'd506  : out_data_ref <= 8'hbb;
      11'd507  : out_data_ref <= 8'h40;
      11'd508  : out_data_ref <= 8'h67;
      11'd509  : out_data_ref <= 8'h90;
      11'd510  : out_data_ref <= 8'h35;
      11'd511  : out_data_ref <= 8'he6;
      11'd512  : out_data_ref <= 8'h52;
      11'd513  : out_data_ref <= 8'h0e;
      11'd514  : out_data_ref <= 8'h09;
      11'd515  : out_data_ref <= 8'hdb;
      11'd516  : out_data_ref <= 8'h91;
      11'd517  : out_data_ref <= 8'hc2;
      11'd518  : out_data_ref <= 8'hf4;
      11'd519  : out_data_ref <= 8'h42;
      11'd520  : out_data_ref <= 8'h72;
      11'd521  : out_data_ref <= 8'h65;
      11'd522  : out_data_ref <= 8'h80;
      11'd523  : out_data_ref <= 8'h6a;
      11'd524  : out_data_ref <= 8'h31;
      11'd525  : out_data_ref <= 8'h41;
      11'd526  : out_data_ref <= 8'h47;
      11'd527  : out_data_ref <= 8'h68;
      11'd528  : out_data_ref <= 8'h74;
      11'd529  : out_data_ref <= 8'h2f;
      11'd530  : out_data_ref <= 8'h34;
      11'd531  : out_data_ref <= 8'h38;
      11'd532  : out_data_ref <= 8'h1c;
      11'd533  : out_data_ref <= 8'h78;
      11'd534  : out_data_ref <= 8'heb;
      11'd535  : out_data_ref <= 8'h9e;
      11'd536  : out_data_ref <= 8'hc7;
      11'd537  : out_data_ref <= 8'ha2;
      11'd538  : out_data_ref <= 8'hbb;
      11'd539  : out_data_ref <= 8'hd3;
      11'd540  : out_data_ref <= 8'ha7;
      11'd541  : out_data_ref <= 8'h03;
      11'd542  : out_data_ref <= 8'hd1;
      11'd543  : out_data_ref <= 8'h3c;
      11'd544  : out_data_ref <= 8'h82;
      11'd545  : out_data_ref <= 8'h90;
      11'd546  : out_data_ref <= 8'hdf;
      11'd547  : out_data_ref <= 8'hf6;
      11'd548  : out_data_ref <= 8'h56;
      11'd549  : out_data_ref <= 8'h69;
      11'd550  : out_data_ref <= 8'h4c;
      11'd551  : out_data_ref <= 8'h32;
      11'd552  : out_data_ref <= 8'h51;
      11'd553  : out_data_ref <= 8'h11;
      11'd554  : out_data_ref <= 8'hef;
      11'd555  : out_data_ref <= 8'h2b;
      11'd556  : out_data_ref <= 8'hed;
      11'd557  : out_data_ref <= 8'h5f;
      11'd558  : out_data_ref <= 8'hd2;
      11'd559  : out_data_ref <= 8'h91;
      11'd560  : out_data_ref <= 8'h32;
      11'd561  : out_data_ref <= 8'h22;
      11'd562  : out_data_ref <= 8'h17;
      11'd563  : out_data_ref <= 8'ha4;
      11'd564  : out_data_ref <= 8'hf9;
      11'd565  : out_data_ref <= 8'h29;
      11'd566  : out_data_ref <= 8'h17;
      11'd567  : out_data_ref <= 8'hcd;
      11'd568  : out_data_ref <= 8'h5d;
      11'd569  : out_data_ref <= 8'h96;
      11'd570  : out_data_ref <= 8'h86;
      11'd571  : out_data_ref <= 8'h75;
      11'd572  : out_data_ref <= 8'he4;
      11'd573  : out_data_ref <= 8'hcb;
      11'd574  : out_data_ref <= 8'hf2;
      11'd575  : out_data_ref <= 8'he8;
      11'd576  : out_data_ref <= 8'h77;
      11'd577  : out_data_ref <= 8'hb7;
      11'd578  : out_data_ref <= 8'he3;
      11'd579  : out_data_ref <= 8'he0;
      11'd580  : out_data_ref <= 8'hbf;
      11'd581  : out_data_ref <= 8'h75;
      11'd582  : out_data_ref <= 8'h94;
      11'd583  : out_data_ref <= 8'h67;
      11'd584  : out_data_ref <= 8'hd1;
      11'd585  : out_data_ref <= 8'hf6;
      11'd586  : out_data_ref <= 8'h98;
      11'd587  : out_data_ref <= 8'h64;
      11'd588  : out_data_ref <= 8'haa;
      11'd589  : out_data_ref <= 8'h1e;
      11'd590  : out_data_ref <= 8'h44;
      11'd591  : out_data_ref <= 8'hcc;
      11'd592  : out_data_ref <= 8'h60;
      11'd593  : out_data_ref <= 8'heb;
      11'd594  : out_data_ref <= 8'hfa;
      11'd595  : out_data_ref <= 8'h2b;
      11'd596  : out_data_ref <= 8'hcf;
      11'd597  : out_data_ref <= 8'h24;
      11'd598  : out_data_ref <= 8'h32;
      11'd599  : out_data_ref <= 8'hfb;
      11'd600  : out_data_ref <= 8'h3b;
      11'd601  : out_data_ref <= 8'h0f;
      11'd602  : out_data_ref <= 8'h09;
      11'd603  : out_data_ref <= 8'h74;
      11'd604  : out_data_ref <= 8'h86;
      11'd605  : out_data_ref <= 8'hb8;
      11'd606  : out_data_ref <= 8'hbd;
      11'd607  : out_data_ref <= 8'hbf;
      11'd608  : out_data_ref <= 8'h0f;
      11'd609  : out_data_ref <= 8'ha9;
      11'd610  : out_data_ref <= 8'h99;
      11'd611  : out_data_ref <= 8'ha4;
      11'd612  : out_data_ref <= 8'he8;
      11'd613  : out_data_ref <= 8'h90;
      11'd614  : out_data_ref <= 8'ha0;
      11'd615  : out_data_ref <= 8'h3b;
      11'd616  : out_data_ref <= 8'h43;
      11'd617  : out_data_ref <= 8'hd8;
      11'd618  : out_data_ref <= 8'h78;
      11'd619  : out_data_ref <= 8'hdd;
      11'd620  : out_data_ref <= 8'hcc;
      11'd621  : out_data_ref <= 8'h3f;
      11'd622  : out_data_ref <= 8'hf0;
      11'd623  : out_data_ref <= 8'h61;
      11'd624  : out_data_ref <= 8'h7a;
      11'd625  : out_data_ref <= 8'h60;
      11'd626  : out_data_ref <= 8'hf8;
      11'd627  : out_data_ref <= 8'h7d;
      11'd628  : out_data_ref <= 8'h49;
      11'd629  : out_data_ref <= 8'h2c;
      11'd630  : out_data_ref <= 8'h10;
      11'd631  : out_data_ref <= 8'h7f;
      11'd632  : out_data_ref <= 8'hdf;
      11'd633  : out_data_ref <= 8'h9e;
      11'd634  : out_data_ref <= 8'h6c;
      11'd635  : out_data_ref <= 8'h86;
      11'd636  : out_data_ref <= 8'hf4;
      11'd637  : out_data_ref <= 8'h76;
      11'd638  : out_data_ref <= 8'hce;
      11'd639  : out_data_ref <= 8'hf9;
      11'd640  : out_data_ref <= 8'hca;
      11'd641  : out_data_ref <= 8'hbe;
      11'd642  : out_data_ref <= 8'hcb;
      11'd643  : out_data_ref <= 8'h6a;
      11'd644  : out_data_ref <= 8'h9c;
      11'd645  : out_data_ref <= 8'h58;
      11'd646  : out_data_ref <= 8'h10;
      11'd647  : out_data_ref <= 8'hab;
      11'd648  : out_data_ref <= 8'h93;
      11'd649  : out_data_ref <= 8'h19;
      11'd650  : out_data_ref <= 8'h8d;
      11'd651  : out_data_ref <= 8'hc8;
      11'd652  : out_data_ref <= 8'h6e;
      11'd653  : out_data_ref <= 8'hef;
      11'd654  : out_data_ref <= 8'he8;
      11'd655  : out_data_ref <= 8'h01;
      11'd656  : out_data_ref <= 8'h51;
      11'd657  : out_data_ref <= 8'h5d;
      11'd658  : out_data_ref <= 8'hb8;
      11'd659  : out_data_ref <= 8'hce;
      11'd660  : out_data_ref <= 8'h96;
      11'd661  : out_data_ref <= 8'ha3;
      11'd662  : out_data_ref <= 8'ha8;
      11'd663  : out_data_ref <= 8'h27;
      11'd664  : out_data_ref <= 8'h0d;
      11'd665  : out_data_ref <= 8'h76;
      11'd666  : out_data_ref <= 8'h1d;
      11'd667  : out_data_ref <= 8'h8b;
      11'd668  : out_data_ref <= 8'h6b;
      11'd669  : out_data_ref <= 8'h94;
      11'd670  : out_data_ref <= 8'h1e;
      11'd671  : out_data_ref <= 8'hd0;
      11'd672  : out_data_ref <= 8'h99;
      11'd673  : out_data_ref <= 8'h9d;
      11'd674  : out_data_ref <= 8'h1e;
      11'd675  : out_data_ref <= 8'h4e;
      11'd676  : out_data_ref <= 8'h65;
      11'd677  : out_data_ref <= 8'hb7;
      11'd678  : out_data_ref <= 8'h4f;
      11'd679  : out_data_ref <= 8'h91;
      11'd680  : out_data_ref <= 8'hee;
      11'd681  : out_data_ref <= 8'h94;
      11'd682  : out_data_ref <= 8'he1;
      11'd683  : out_data_ref <= 8'hc9;
      11'd684  : out_data_ref <= 8'h90;
      11'd685  : out_data_ref <= 8'h38;
      11'd686  : out_data_ref <= 8'hd6;
      11'd687  : out_data_ref <= 8'hbf;
      11'd688  : out_data_ref <= 8'he7;
      11'd689  : out_data_ref <= 8'hd6;
      11'd690  : out_data_ref <= 8'h24;
      11'd691  : out_data_ref <= 8'hcc;
      11'd692  : out_data_ref <= 8'h64;
      11'd693  : out_data_ref <= 8'h7a;
      11'd694  : out_data_ref <= 8'hbd;
      11'd695  : out_data_ref <= 8'h84;
      11'd696  : out_data_ref <= 8'h54;
      11'd697  : out_data_ref <= 8'h18;
      11'd698  : out_data_ref <= 8'h5d;
      11'd699  : out_data_ref <= 8'h8a;
      11'd700  : out_data_ref <= 8'h89;
      11'd701  : out_data_ref <= 8'hb2;
      11'd702  : out_data_ref <= 8'h58;
      11'd703  : out_data_ref <= 8'h1b;
      11'd704  : out_data_ref <= 8'h82;
      11'd705  : out_data_ref <= 8'he1;
      11'd706  : out_data_ref <= 8'h88;
      11'd707  : out_data_ref <= 8'h63;
      11'd708  : out_data_ref <= 8'h36;
      11'd709  : out_data_ref <= 8'hcb;
      11'd710  : out_data_ref <= 8'h47;
      11'd711  : out_data_ref <= 8'h36;
      11'd712  : out_data_ref <= 8'h89;
      11'd713  : out_data_ref <= 8'hda;
      11'd714  : out_data_ref <= 8'h83;
      11'd715  : out_data_ref <= 8'h38;
      11'd716  : out_data_ref <= 8'h64;
      11'd717  : out_data_ref <= 8'he5;
      11'd718  : out_data_ref <= 8'h27;
      11'd719  : out_data_ref <= 8'h98;
      11'd720  : out_data_ref <= 8'h17;
      11'd721  : out_data_ref <= 8'hf1;
      11'd722  : out_data_ref <= 8'h41;
      11'd723  : out_data_ref <= 8'h1c;
      11'd724  : out_data_ref <= 8'hb8;
      11'd725  : out_data_ref <= 8'he1;
      11'd726  : out_data_ref <= 8'h1d;
      11'd727  : out_data_ref <= 8'h9a;
      11'd728  : out_data_ref <= 8'h20;
      11'd729  : out_data_ref <= 8'h1e;
      11'd730  : out_data_ref <= 8'hee;
      11'd731  : out_data_ref <= 8'h51;
      11'd732  : out_data_ref <= 8'h33;
      11'd733  : out_data_ref <= 8'he2;
      11'd734  : out_data_ref <= 8'h70;
      11'd735  : out_data_ref <= 8'hf4;
      11'd736  : out_data_ref <= 8'h99;
      11'd737  : out_data_ref <= 8'h1e;
      11'd738  : out_data_ref <= 8'hbd;
      11'd739  : out_data_ref <= 8'h17;
      11'd740  : out_data_ref <= 8'h9f;
      11'd741  : out_data_ref <= 8'h5d;
      11'd742  : out_data_ref <= 8'ha0;
      11'd743  : out_data_ref <= 8'h0b;
      11'd744  : out_data_ref <= 8'h2e;
      11'd745  : out_data_ref <= 8'h73;
      11'd746  : out_data_ref <= 8'h3d;
      11'd747  : out_data_ref <= 8'h59;
      11'd748  : out_data_ref <= 8'hc8;
      11'd749  : out_data_ref <= 8'hab;
      11'd750  : out_data_ref <= 8'h65;
      11'd751  : out_data_ref <= 8'h6c;
      11'd752  : out_data_ref <= 8'h40;
      11'd753  : out_data_ref <= 8'h2f;
      11'd754  : out_data_ref <= 8'he0;
      11'd755  : out_data_ref <= 8'hdd;
      11'd756  : out_data_ref <= 8'ha2;
      11'd757  : out_data_ref <= 8'h1c;
      11'd758  : out_data_ref <= 8'h97;
      11'd759  : out_data_ref <= 8'heb;
      11'd760  : out_data_ref <= 8'ha1;
      11'd761  : out_data_ref <= 8'hfc;
      11'd762  : out_data_ref <= 8'hc4;
      11'd763  : out_data_ref <= 8'h16;
      11'd764  : out_data_ref <= 8'h1e;
      11'd765  : out_data_ref <= 8'h49;
      11'd766  : out_data_ref <= 8'hb1;
      11'd767  : out_data_ref <= 8'ha4;
      11'd768  : out_data_ref <= 8'h55;
      11'd769  : out_data_ref <= 8'h74;
      11'd770  : out_data_ref <= 8'h75;
      11'd771  : out_data_ref <= 8'h0b;
      11'd772  : out_data_ref <= 8'h5f;
      11'd773  : out_data_ref <= 8'h00;
      11'd774  : out_data_ref <= 8'h78;
      11'd775  : out_data_ref <= 8'h23;
      11'd776  : out_data_ref <= 8'h42;
      11'd777  : out_data_ref <= 8'hae;
      11'd778  : out_data_ref <= 8'hc2;
      11'd779  : out_data_ref <= 8'h2a;
      11'd780  : out_data_ref <= 8'h08;
      11'd781  : out_data_ref <= 8'hb4;
      11'd782  : out_data_ref <= 8'haa;
      11'd783  : out_data_ref <= 8'h4a;
      11'd784  : out_data_ref <= 8'h73;
      11'd785  : out_data_ref <= 8'he7;
      11'd786  : out_data_ref <= 8'h57;
      11'd787  : out_data_ref <= 8'h2e;
      11'd788  : out_data_ref <= 8'h3a;
      11'd789  : out_data_ref <= 8'hcd;
      11'd790  : out_data_ref <= 8'h95;
      11'd791  : out_data_ref <= 8'h9c;
      11'd792  : out_data_ref <= 8'h4a;
      11'd793  : out_data_ref <= 8'hd2;
      11'd794  : out_data_ref <= 8'hd5;
      11'd795  : out_data_ref <= 8'h50;
      11'd796  : out_data_ref <= 8'h1b;
      11'd797  : out_data_ref <= 8'hc0;
      11'd798  : out_data_ref <= 8'ha6;
      11'd799  : out_data_ref <= 8'h02;
      11'd800  : out_data_ref <= 8'h7b;
      11'd801  : out_data_ref <= 8'hdc;
      11'd802  : out_data_ref <= 8'h09;
      11'd803  : out_data_ref <= 8'h1c;
      11'd804  : out_data_ref <= 8'hb1;
      11'd805  : out_data_ref <= 8'h08;
      11'd806  : out_data_ref <= 8'hcc;
      11'd807  : out_data_ref <= 8'h99;
      11'd808  : out_data_ref <= 8'h4f;
      11'd809  : out_data_ref <= 8'hcf;
      11'd810  : out_data_ref <= 8'he4;
      11'd811  : out_data_ref <= 8'h8c;
      11'd812  : out_data_ref <= 8'hcc;
      11'd813  : out_data_ref <= 8'h89;
      11'd814  : out_data_ref <= 8'h6f;
      11'd815  : out_data_ref <= 8'h21;
      11'd816  : out_data_ref <= 8'h52;
      11'd817  : out_data_ref <= 8'h5e;
      11'd818  : out_data_ref <= 8'h89;
      11'd819  : out_data_ref <= 8'h85;
      11'd820  : out_data_ref <= 8'hfc;
      11'd821  : out_data_ref <= 8'had;
      11'd822  : out_data_ref <= 8'hc8;
      11'd823  : out_data_ref <= 8'h12;
      11'd824  : out_data_ref <= 8'h69;
      11'd825  : out_data_ref <= 8'h40;
      11'd826  : out_data_ref <= 8'he3;
      11'd827  : out_data_ref <= 8'hd4;
      11'd828  : out_data_ref <= 8'h57;
      11'd829  : out_data_ref <= 8'h6b;
      11'd830  : out_data_ref <= 8'hb5;
      11'd831  : out_data_ref <= 8'hb4;
      11'd832  : out_data_ref <= 8'hfd;
      11'd833  : out_data_ref <= 8'hc6;
      11'd834  : out_data_ref <= 8'h08;
      11'd835  : out_data_ref <= 8'h6a;
      11'd836  : out_data_ref <= 8'hc0;
      11'd837  : out_data_ref <= 8'he9;
      11'd838  : out_data_ref <= 8'he5;
      11'd839  : out_data_ref <= 8'h86;
      11'd840  : out_data_ref <= 8'he9;
      11'd841  : out_data_ref <= 8'hb0;
      11'd842  : out_data_ref <= 8'h55;
      11'd843  : out_data_ref <= 8'ha3;
      11'd844  : out_data_ref <= 8'ha7;
      11'd845  : out_data_ref <= 8'h81;
      11'd846  : out_data_ref <= 8'h0d;
      11'd847  : out_data_ref <= 8'h12;
      11'd848  : out_data_ref <= 8'h17;
      11'd849  : out_data_ref <= 8'h10;
      11'd850  : out_data_ref <= 8'hcf;
      11'd851  : out_data_ref <= 8'h8c;
      11'd852  : out_data_ref <= 8'hf5;
      11'd853  : out_data_ref <= 8'h52;
      11'd854  : out_data_ref <= 8'h3c;
      11'd855  : out_data_ref <= 8'hc4;
      11'd856  : out_data_ref <= 8'h61;
      11'd857  : out_data_ref <= 8'h37;
      11'd858  : out_data_ref <= 8'h55;
      11'd859  : out_data_ref <= 8'hc4;
      11'd860  : out_data_ref <= 8'h9b;
      11'd861  : out_data_ref <= 8'h00;
      11'd862  : out_data_ref <= 8'hef;
      11'd863  : out_data_ref <= 8'h36;
      11'd864  : out_data_ref <= 8'hc1;
      11'd865  : out_data_ref <= 8'h61;
      11'd866  : out_data_ref <= 8'h2c;
      11'd867  : out_data_ref <= 8'h0f;
      11'd868  : out_data_ref <= 8'hae;
      11'd869  : out_data_ref <= 8'hda;
      11'd870  : out_data_ref <= 8'hac;
      11'd871  : out_data_ref <= 8'h31;
      11'd872  : out_data_ref <= 8'h39;
      11'd873  : out_data_ref <= 8'h63;
      11'd874  : out_data_ref <= 8'hdd;
      11'd875  : out_data_ref <= 8'h34;
      11'd876  : out_data_ref <= 8'h55;
      11'd877  : out_data_ref <= 8'hfc;
      11'd878  : out_data_ref <= 8'h9f;
      11'd879  : out_data_ref <= 8'h81;
      11'd880  : out_data_ref <= 8'h34;
      11'd881  : out_data_ref <= 8'hb8;
      11'd882  : out_data_ref <= 8'h4b;
      11'd883  : out_data_ref <= 8'hd0;
      11'd884  : out_data_ref <= 8'hb8;
      11'd885  : out_data_ref <= 8'h02;
      11'd886  : out_data_ref <= 8'h12;
      11'd887  : out_data_ref <= 8'h5d;
      11'd888  : out_data_ref <= 8'h4c;
      11'd889  : out_data_ref <= 8'h20;
      11'd890  : out_data_ref <= 8'h12;
      11'd891  : out_data_ref <= 8'h6f;
      11'd892  : out_data_ref <= 8'hbe;
      11'd893  : out_data_ref <= 8'hd4;
      11'd894  : out_data_ref <= 8'hf7;
      11'd895  : out_data_ref <= 8'h30;
      11'd896  : out_data_ref <= 8'h13;
      11'd897  : out_data_ref <= 8'h95;
      11'd898  : out_data_ref <= 8'h38;
      11'd899  : out_data_ref <= 8'hd6;
      11'd900  : out_data_ref <= 8'hc3;
      11'd901  : out_data_ref <= 8'h6b;
      11'd902  : out_data_ref <= 8'hc4;
      11'd903  : out_data_ref <= 8'h0e;
      11'd904  : out_data_ref <= 8'hde;
      11'd905  : out_data_ref <= 8'hdf;
      11'd906  : out_data_ref <= 8'h0b;
      11'd907  : out_data_ref <= 8'h8d;
      11'd908  : out_data_ref <= 8'hbb;
      11'd909  : out_data_ref <= 8'h8c;
      11'd910  : out_data_ref <= 8'hd3;
      11'd911  : out_data_ref <= 8'h15;
      11'd912  : out_data_ref <= 8'h00;
      11'd913  : out_data_ref <= 8'h03;
      11'd914  : out_data_ref <= 8'hb2;
      11'd915  : out_data_ref <= 8'h8e;
      11'd916  : out_data_ref <= 8'h2d;
      11'd917  : out_data_ref <= 8'h32;
      11'd918  : out_data_ref <= 8'ha3;
      11'd919  : out_data_ref <= 8'h77;
      11'd920  : out_data_ref <= 8'hb3;
      11'd921  : out_data_ref <= 8'hb8;
      11'd922  : out_data_ref <= 8'h99;
      11'd923  : out_data_ref <= 8'hb2;
      11'd924  : out_data_ref <= 8'ha1;
      11'd925  : out_data_ref <= 8'h93;
      11'd926  : out_data_ref <= 8'hcb;
      11'd927  : out_data_ref <= 8'he0;
      11'd928  : out_data_ref <= 8'h5f;
      11'd929  : out_data_ref <= 8'hfa;
      11'd930  : out_data_ref <= 8'h57;
      11'd931  : out_data_ref <= 8'h6a;
      11'd932  : out_data_ref <= 8'h2c;
      11'd933  : out_data_ref <= 8'h48;
      11'd934  : out_data_ref <= 8'he5;
      11'd935  : out_data_ref <= 8'hdc;
      11'd936  : out_data_ref <= 8'h76;
      11'd937  : out_data_ref <= 8'hb8;
      11'd938  : out_data_ref <= 8'h4e;
      11'd939  : out_data_ref <= 8'h89;
      11'd940  : out_data_ref <= 8'hcf;
      11'd941  : out_data_ref <= 8'h87;
      11'd942  : out_data_ref <= 8'hb3;
      11'd943  : out_data_ref <= 8'hee;
      11'd944  : out_data_ref <= 8'he0;
      11'd945  : out_data_ref <= 8'h56;
      11'd946  : out_data_ref <= 8'h3b;
      11'd947  : out_data_ref <= 8'h47;
      11'd948  : out_data_ref <= 8'h7e;
      11'd949  : out_data_ref <= 8'h0a;
      11'd950  : out_data_ref <= 8'h07;
      11'd951  : out_data_ref <= 8'hdf;
      11'd952  : out_data_ref <= 8'h43;
      11'd953  : out_data_ref <= 8'h3f;
      11'd954  : out_data_ref <= 8'h4e;
      11'd955  : out_data_ref <= 8'hec;
      11'd956  : out_data_ref <= 8'h3b;
      11'd957  : out_data_ref <= 8'h20;
      11'd958  : out_data_ref <= 8'hf0;
      11'd959  : out_data_ref <= 8'hb0;
      11'd960  : out_data_ref <= 8'h12;
      11'd961  : out_data_ref <= 8'hf4;
      11'd962  : out_data_ref <= 8'hb5;
      11'd963  : out_data_ref <= 8'hae;
      11'd964  : out_data_ref <= 8'h11;
      11'd965  : out_data_ref <= 8'h1c;
      11'd966  : out_data_ref <= 8'h2f;
      11'd967  : out_data_ref <= 8'hf6;
      11'd968  : out_data_ref <= 8'hee;
      11'd969  : out_data_ref <= 8'h5b;
      11'd970  : out_data_ref <= 8'hcd;
      11'd971  : out_data_ref <= 8'he9;
      11'd972  : out_data_ref <= 8'ha3;
      11'd973  : out_data_ref <= 8'he5;
      11'd974  : out_data_ref <= 8'hfc;
      11'd975  : out_data_ref <= 8'hbb;
      11'd976  : out_data_ref <= 8'h76;
      11'd977  : out_data_ref <= 8'h7c;
      11'd978  : out_data_ref <= 8'hfa;
      11'd979  : out_data_ref <= 8'h4f;
      11'd980  : out_data_ref <= 8'hb8;
      11'd981  : out_data_ref <= 8'ha3;
      11'd982  : out_data_ref <= 8'hdb;
      11'd983  : out_data_ref <= 8'hc8;
      11'd984  : out_data_ref <= 8'hf5;
      11'd985  : out_data_ref <= 8'h6a;
      11'd986  : out_data_ref <= 8'h46;
      11'd987  : out_data_ref <= 8'h81;
      11'd988  : out_data_ref <= 8'h77;
      11'd989  : out_data_ref <= 8'hf2;
      11'd990  : out_data_ref <= 8'heb;
      11'd991  : out_data_ref <= 8'h2a;
      11'd992  : out_data_ref <= 8'hd2;
      11'd993  : out_data_ref <= 8'h72;
      11'd994  : out_data_ref <= 8'h0c;
      11'd995  : out_data_ref <= 8'h7c;
      11'd996  : out_data_ref <= 8'hfb;
      11'd997  : out_data_ref <= 8'h83;
      11'd998  : out_data_ref <= 8'hb5;
      11'd999  : out_data_ref <= 8'hda;
      11'd1000 : out_data_ref <= 8'h90;
      11'd1001 : out_data_ref <= 8'h4a;
      11'd1002 : out_data_ref <= 8'hbb;
      11'd1003 : out_data_ref <= 8'hd6;
      11'd1004 : out_data_ref <= 8'hbb;
      11'd1005 : out_data_ref <= 8'h67;
      11'd1006 : out_data_ref <= 8'h1a;
      11'd1007 : out_data_ref <= 8'hf8;
      11'd1008 : out_data_ref <= 8'hc3;
      11'd1009 : out_data_ref <= 8'h33;
      11'd1010 : out_data_ref <= 8'ha2;
      11'd1011 : out_data_ref <= 8'hef;
      11'd1012 : out_data_ref <= 8'h9a;
      11'd1013 : out_data_ref <= 8'h8b;
      11'd1014 : out_data_ref <= 8'hf5;
      11'd1015 : out_data_ref <= 8'h6f;
      11'd1016 : out_data_ref <= 8'hb8;
      11'd1017 : out_data_ref <= 8'h0c;
      11'd1018 : out_data_ref <= 8'h9b;
      11'd1019 : out_data_ref <= 8'hd7;
      11'd1020 : out_data_ref <= 8'h99;
      11'd1021 : out_data_ref <= 8'hff;
      11'd1022 : out_data_ref <= 8'hf4;
      11'd1023 : out_data_ref <= 8'h58;
      11'd1024 : out_data_ref <= 8'h6e;
      11'd1025 : out_data_ref <= 8'h65;
      11'd1026 : out_data_ref <= 8'h68;
      11'd1027 : out_data_ref <= 8'h16;
      11'd1028 : out_data_ref <= 8'hbb;
      11'd1029 : out_data_ref <= 8'h76;
      11'd1030 : out_data_ref <= 8'hdb;
      11'd1031 : out_data_ref <= 8'hb7;
      11'd1032 : out_data_ref <= 8'ha7;
      11'd1033 : out_data_ref <= 8'hd8;
      11'd1034 : out_data_ref <= 8'h0e;
      11'd1035 : out_data_ref <= 8'h70;
      11'd1036 : out_data_ref <= 8'h01;
      11'd1037 : out_data_ref <= 8'hb5;
      11'd1038 : out_data_ref <= 8'he5;
      11'd1039 : out_data_ref <= 8'h99;
      11'd1040 : out_data_ref <= 8'ha5;
      11'd1041 : out_data_ref <= 8'h62;
      11'd1042 : out_data_ref <= 8'ha3;
      11'd1043 : out_data_ref <= 8'h64;
      11'd1044 : out_data_ref <= 8'ha5;
      11'd1045 : out_data_ref <= 8'h0c;
      11'd1046 : out_data_ref <= 8'h5e;
      11'd1047 : out_data_ref <= 8'h89;
      11'd1048 : out_data_ref <= 8'h49;
      11'd1049 : out_data_ref <= 8'hfa;
      11'd1050 : out_data_ref <= 8'h5a;
      11'd1051 : out_data_ref <= 8'h18;
      11'd1052 : out_data_ref <= 8'h4d;
      11'd1053 : out_data_ref <= 8'h8e;
      11'd1054 : out_data_ref <= 8'had;
      11'd1055 : out_data_ref <= 8'h72;
      11'd1056 : out_data_ref <= 8'hf2;
      11'd1057 : out_data_ref <= 8'h98;
      11'd1058 : out_data_ref <= 8'hdd;
      11'd1059 : out_data_ref <= 8'h7c;
      11'd1060 : out_data_ref <= 8'h84;
      11'd1061 : out_data_ref <= 8'h13;
      11'd1062 : out_data_ref <= 8'h07;
      11'd1063 : out_data_ref <= 8'h1c;
      11'd1064 : out_data_ref <= 8'h51;
      11'd1065 : out_data_ref <= 8'hed;
      11'd1066 : out_data_ref <= 8'had;
      11'd1067 : out_data_ref <= 8'hc8;
      11'd1068 : out_data_ref <= 8'h18;
      11'd1069 : out_data_ref <= 8'h53;
      11'd1070 : out_data_ref <= 8'ha7;
      11'd1071 : out_data_ref <= 8'h40;
      11'd1072 : out_data_ref <= 8'h04;
      11'd1073 : out_data_ref <= 8'hcc;
      11'd1074 : out_data_ref <= 8'ha6;
      11'd1075 : out_data_ref <= 8'h89;
      11'd1076 : out_data_ref <= 8'h1b;
      11'd1077 : out_data_ref <= 8'hbd;
      11'd1078 : out_data_ref <= 8'h10;
      11'd1079 : out_data_ref <= 8'h1c;
      11'd1080 : out_data_ref <= 8'h6b;
      11'd1081 : out_data_ref <= 8'h65;
      11'd1082 : out_data_ref <= 8'haf;
      11'd1083 : out_data_ref <= 8'h35;
      11'd1084 : out_data_ref <= 8'ha6;
      11'd1085 : out_data_ref <= 8'h2a;
      11'd1086 : out_data_ref <= 8'h5b;
      11'd1087 : out_data_ref <= 8'h2b;
      11'd1088 : out_data_ref <= 8'hf5;
      11'd1089 : out_data_ref <= 8'h43;
      11'd1090 : out_data_ref <= 8'h06;
      11'd1091 : out_data_ref <= 8'he1;
      11'd1092 : out_data_ref <= 8'h8d;
      11'd1093 : out_data_ref <= 8'h10;
      11'd1094 : out_data_ref <= 8'h16;
      11'd1095 : out_data_ref <= 8'h8a;
      11'd1096 : out_data_ref <= 8'hc8;
      11'd1097 : out_data_ref <= 8'h9d;
      11'd1098 : out_data_ref <= 8'h93;
      11'd1099 : out_data_ref <= 8'h6e;
      11'd1100 : out_data_ref <= 8'h03;
      11'd1101 : out_data_ref <= 8'h85;
      11'd1102 : out_data_ref <= 8'h0d;
      11'd1103 : out_data_ref <= 8'h89;
      11'd1104 : out_data_ref <= 8'h94;
      11'd1105 : out_data_ref <= 8'h1e;
      11'd1106 : out_data_ref <= 8'h60;
      11'd1107 : out_data_ref <= 8'hd1;
      11'd1108 : out_data_ref <= 8'hf4;
      11'd1109 : out_data_ref <= 8'h4b;
      11'd1110 : out_data_ref <= 8'h02;
      11'd1111 : out_data_ref <= 8'h0b;
      11'd1112 : out_data_ref <= 8'h87;
      11'd1113 : out_data_ref <= 8'he1;
      11'd1114 : out_data_ref <= 8'h5f;
      11'd1115 : out_data_ref <= 8'h77;
      11'd1116 : out_data_ref <= 8'hec;
      11'd1117 : out_data_ref <= 8'h6d;
      11'd1118 : out_data_ref <= 8'h6c;
      11'd1119 : out_data_ref <= 8'h0e;
      11'd1120 : out_data_ref <= 8'h4b;
      11'd1121 : out_data_ref <= 8'hef;
      11'd1122 : out_data_ref <= 8'h99;
      11'd1123 : out_data_ref <= 8'h70;
      11'd1124 : out_data_ref <= 8'h57;
      11'd1125 : out_data_ref <= 8'h9b;
      11'd1126 : out_data_ref <= 8'h15;
      11'd1127 : out_data_ref <= 8'h38;
      11'd1128 : out_data_ref <= 8'h88;
      11'd1129 : out_data_ref <= 8'h64;
      11'd1130 : out_data_ref <= 8'h66;
      11'd1131 : out_data_ref <= 8'hb1;
      11'd1132 : out_data_ref <= 8'h79;
      11'd1133 : out_data_ref <= 8'h43;
      11'd1134 : out_data_ref <= 8'ha8;
      11'd1135 : out_data_ref <= 8'h9c;
      11'd1136 : out_data_ref <= 8'h23;
      11'd1137 : out_data_ref <= 8'h39;
      11'd1138 : out_data_ref <= 8'hc9;
      11'd1139 : out_data_ref <= 8'h7f;
      11'd1140 : out_data_ref <= 8'h6d;
      11'd1141 : out_data_ref <= 8'h65;
      11'd1142 : out_data_ref <= 8'h69;
      11'd1143 : out_data_ref <= 8'h5a;
      11'd1144 : out_data_ref <= 8'h4d;
      11'd1145 : out_data_ref <= 8'h3d;
      11'd1146 : out_data_ref <= 8'he3;
      11'd1147 : out_data_ref <= 8'h64;
      11'd1148 : out_data_ref <= 8'ha4;
      11'd1149 : out_data_ref <= 8'hd1;
      11'd1150 : out_data_ref <= 8'hb0;
      11'd1151 : out_data_ref <= 8'hbe;
      11'd1152 : out_data_ref <= 8'h80;
      11'd1153 : out_data_ref <= 8'h10;
      11'd1154 : out_data_ref <= 8'h87;
      11'd1155 : out_data_ref <= 8'h6d;
      11'd1156 : out_data_ref <= 8'h67;
      11'd1157 : out_data_ref <= 8'he3;
      11'd1158 : out_data_ref <= 8'h1c;
      11'd1159 : out_data_ref <= 8'hb1;
      11'd1160 : out_data_ref <= 8'h1d;
      11'd1161 : out_data_ref <= 8'h67;
      11'd1162 : out_data_ref <= 8'h27;
      11'd1163 : out_data_ref <= 8'h3a;
      11'd1164 : out_data_ref <= 8'hf9;
      11'd1165 : out_data_ref <= 8'hdc;
      11'd1166 : out_data_ref <= 8'h91;
      11'd1167 : out_data_ref <= 8'hfd;
      11'd1168 : out_data_ref <= 8'h19;
      11'd1169 : out_data_ref <= 8'hbe;
      11'd1170 : out_data_ref <= 8'h63;
      11'd1171 : out_data_ref <= 8'h4f;
      11'd1172 : out_data_ref <= 8'h1f;
      11'd1173 : out_data_ref <= 8'hf4;
      11'd1174 : out_data_ref <= 8'hd0;
      11'd1175 : out_data_ref <= 8'hc6;
      11'd1176 : out_data_ref <= 8'h6f;
      11'd1177 : out_data_ref <= 8'h3f;
      11'd1178 : out_data_ref <= 8'h6d;
      11'd1179 : out_data_ref <= 8'h88;
      11'd1180 : out_data_ref <= 8'h2e;
      11'd1181 : out_data_ref <= 8'h51;
      11'd1182 : out_data_ref <= 8'h44;
      11'd1183 : out_data_ref <= 8'h68;
      11'd1184 : out_data_ref <= 8'h8c;
      11'd1185 : out_data_ref <= 8'h27;
      11'd1186 : out_data_ref <= 8'h6b;
      11'd1187 : out_data_ref <= 8'h36;
      11'd1188 : out_data_ref <= 8'h4e;
      11'd1189 : out_data_ref <= 8'h44;
      11'd1190 : out_data_ref <= 8'hd3;
      11'd1191 : out_data_ref <= 8'hb3;
      11'd1192 : out_data_ref <= 8'h8c;
      11'd1193 : out_data_ref <= 8'hd2;
      11'd1194 : out_data_ref <= 8'h62;
      11'd1195 : out_data_ref <= 8'h06;
      11'd1196 : out_data_ref <= 8'h42;
      11'd1197 : out_data_ref <= 8'h20;
      11'd1198 : out_data_ref <= 8'hc4;
      11'd1199 : out_data_ref <= 8'h27;
      11'd1200 : out_data_ref <= 8'h89;
      11'd1201 : out_data_ref <= 8'hdc;
      11'd1202 : out_data_ref <= 8'he9;
      11'd1203 : out_data_ref <= 8'h04;
      11'd1204 : out_data_ref <= 8'h42;
      11'd1205 : out_data_ref <= 8'h25;
      11'd1206 : out_data_ref <= 8'h62;
      11'd1207 : out_data_ref <= 8'h1a;
      11'd1208 : out_data_ref <= 8'hf7;
      11'd1209 : out_data_ref <= 8'h43;
      11'd1210 : out_data_ref <= 8'hd9;
      11'd1211 : out_data_ref <= 8'h8a;
      11'd1212 : out_data_ref <= 8'hed;
      11'd1213 : out_data_ref <= 8'haa;
      11'd1214 : out_data_ref <= 8'h6d;
      11'd1215 : out_data_ref <= 8'h8d;
      11'd1216 : out_data_ref <= 8'h0e;
      11'd1217 : out_data_ref <= 8'h59;
      11'd1218 : out_data_ref <= 8'h25;
      11'd1219 : out_data_ref <= 8'h53;
      11'd1220 : out_data_ref <= 8'hab;
      11'd1221 : out_data_ref <= 8'h4d;
      11'd1222 : out_data_ref <= 8'h45;
      11'd1223 : out_data_ref <= 8'h05;
      11'd1224 : out_data_ref <= 8'h11;
      11'd1225 : out_data_ref <= 8'h25;
      11'd1226 : out_data_ref <= 8'h23;
      11'd1227 : out_data_ref <= 8'hb1;
      11'd1228 : out_data_ref <= 8'h29;
      11'd1229 : out_data_ref <= 8'ha1;
      11'd1230 : out_data_ref <= 8'h65;
      11'd1231 : out_data_ref <= 8'h38;
      11'd1232 : out_data_ref <= 8'h6a;
      11'd1233 : out_data_ref <= 8'hbe;
      11'd1234 : out_data_ref <= 8'h81;
      11'd1235 : out_data_ref <= 8'hf0;
      11'd1236 : out_data_ref <= 8'hec;
      11'd1237 : out_data_ref <= 8'h76;
      11'd1238 : out_data_ref <= 8'hf1;
      11'd1239 : out_data_ref <= 8'hd6;
      11'd1240 : out_data_ref <= 8'he8;
      11'd1241 : out_data_ref <= 8'h76;
      11'd1242 : out_data_ref <= 8'h93;
      11'd1243 : out_data_ref <= 8'h55;
      11'd1244 : out_data_ref <= 8'h54;
      11'd1245 : out_data_ref <= 8'h08;
      11'd1246 : out_data_ref <= 8'h4d;
      11'd1247 : out_data_ref <= 8'h62;
      11'd1248 : out_data_ref <= 8'h08;
      11'd1249 : out_data_ref <= 8'h6e;
      11'd1250 : out_data_ref <= 8'h54;
      11'd1251 : out_data_ref <= 8'h07;
      11'd1252 : out_data_ref <= 8'h0e;
      11'd1253 : out_data_ref <= 8'h11;
      11'd1254 : out_data_ref <= 8'h46;
      11'd1255 : out_data_ref <= 8'h64;
      11'd1256 : out_data_ref <= 8'hd0;
      11'd1257 : out_data_ref <= 8'h79;
      11'd1258 : out_data_ref <= 8'h8e;
      11'd1259 : out_data_ref <= 8'h30;
      11'd1260 : out_data_ref <= 8'h36;
      11'd1261 : out_data_ref <= 8'h7e;
      11'd1262 : out_data_ref <= 8'h30;
      11'd1263 : out_data_ref <= 8'hc9;
      11'd1264 : out_data_ref <= 8'h8f;
      11'd1265 : out_data_ref <= 8'h16;
      11'd1266 : out_data_ref <= 8'hb5;
      11'd1267 : out_data_ref <= 8'h14;
      11'd1268 : out_data_ref <= 8'h77;
      11'd1269 : out_data_ref <= 8'hef;
      11'd1270 : out_data_ref <= 8'hb3;
      11'd1271 : out_data_ref <= 8'h17;
      11'd1272 : out_data_ref <= 8'hbe;
      11'd1273 : out_data_ref <= 8'h15;
      11'd1274 : out_data_ref <= 8'h20;
      11'd1275 : out_data_ref <= 8'h94;
      11'd1276 : out_data_ref <= 8'hc9;
      11'd1277 : out_data_ref <= 8'h97;
      11'd1278 : out_data_ref <= 8'hec;
      11'd1279 : out_data_ref <= 8'h8e;
      11'd1280 : out_data_ref <= 8'hfc;
      11'd1281 : out_data_ref <= 8'hac;
      11'd1282 : out_data_ref <= 8'h33;
      11'd1283 : out_data_ref <= 8'hc9;
      11'd1284 : out_data_ref <= 8'h16;
      11'd1285 : out_data_ref <= 8'he4;
      11'd1286 : out_data_ref <= 8'h1f;
      11'd1287 : out_data_ref <= 8'h63;
      11'd1288 : out_data_ref <= 8'hbd;
      11'd1289 : out_data_ref <= 8'h89;
      11'd1290 : out_data_ref <= 8'h9f;
      11'd1291 : out_data_ref <= 8'h92;
      11'd1292 : out_data_ref <= 8'h77;
      11'd1293 : out_data_ref <= 8'hf1;
      11'd1294 : out_data_ref <= 8'h7d;
      11'd1295 : out_data_ref <= 8'hf4;
      11'd1296 : out_data_ref <= 8'h51;
      11'd1297 : out_data_ref <= 8'h88;
      11'd1298 : out_data_ref <= 8'h93;
      11'd1299 : out_data_ref <= 8'h08;
      11'd1300 : out_data_ref <= 8'h6e;
      11'd1301 : out_data_ref <= 8'h60;
      11'd1302 : out_data_ref <= 8'h12;
      11'd1303 : out_data_ref <= 8'h7c;
      11'd1304 : out_data_ref <= 8'hc5;
      11'd1305 : out_data_ref <= 8'hdc;
      11'd1306 : out_data_ref <= 8'h18;
      11'd1307 : out_data_ref <= 8'h31;
      11'd1308 : out_data_ref <= 8'he8;
      11'd1309 : out_data_ref <= 8'h55;
      11'd1310 : out_data_ref <= 8'hb1;
      11'd1311 : out_data_ref <= 8'ha0;
      11'd1312 : out_data_ref <= 8'h82;
      11'd1313 : out_data_ref <= 8'h72;
      11'd1314 : out_data_ref <= 8'hb6;
      11'd1315 : out_data_ref <= 8'had;
      11'd1316 : out_data_ref <= 8'hd9;
      11'd1317 : out_data_ref <= 8'h6d;
      11'd1318 : out_data_ref <= 8'hfc;
      11'd1319 : out_data_ref <= 8'h5d;
      11'd1320 : out_data_ref <= 8'ha0;
      11'd1321 : out_data_ref <= 8'h17;
      11'd1322 : out_data_ref <= 8'he1;
      11'd1323 : out_data_ref <= 8'h78;
      11'd1324 : out_data_ref <= 8'h3a;
      11'd1325 : out_data_ref <= 8'hc0;
      11'd1326 : out_data_ref <= 8'hfd;
      11'd1327 : out_data_ref <= 8'h81;
      11'd1328 : out_data_ref <= 8'h37;
      11'd1329 : out_data_ref <= 8'hfb;
      11'd1330 : out_data_ref <= 8'h65;
      11'd1331 : out_data_ref <= 8'hed;
      11'd1332 : out_data_ref <= 8'hbc;
      11'd1333 : out_data_ref <= 8'hb9;
      11'd1334 : out_data_ref <= 8'h70;
      11'd1335 : out_data_ref <= 8'h0f;
      11'd1336 : out_data_ref <= 8'h04;
      11'd1337 : out_data_ref <= 8'h39;
      11'd1338 : out_data_ref <= 8'hc6;
      11'd1339 : out_data_ref <= 8'hf1;
      11'd1340 : out_data_ref <= 8'h1b;
      11'd1341 : out_data_ref <= 8'hbb;
      11'd1342 : out_data_ref <= 8'h62;
      11'd1343 : out_data_ref <= 8'hc7;
      11'd1344 : out_data_ref <= 8'h36;
      11'd1345 : out_data_ref <= 8'h00;
      11'd1346 : out_data_ref <= 8'h15;
      11'd1347 : out_data_ref <= 8'h98;
      11'd1348 : out_data_ref <= 8'h01;
      11'd1349 : out_data_ref <= 8'hc2;
      11'd1350 : out_data_ref <= 8'had;
      11'd1351 : out_data_ref <= 8'hf2;
      11'd1352 : out_data_ref <= 8'h57;
      11'd1353 : out_data_ref <= 8'hda;
      11'd1354 : out_data_ref <= 8'ha1;
      11'd1355 : out_data_ref <= 8'h92;
      11'd1356 : out_data_ref <= 8'hfe;
      11'd1357 : out_data_ref <= 8'hfc;
      11'd1358 : out_data_ref <= 8'h6a;
      11'd1359 : out_data_ref <= 8'hdf;
      11'd1360 : out_data_ref <= 8'hf9;
      11'd1361 : out_data_ref <= 8'h64;
      11'd1362 : out_data_ref <= 8'h86;
      11'd1363 : out_data_ref <= 8'hd6;
      11'd1364 : out_data_ref <= 8'he6;
      11'd1365 : out_data_ref <= 8'h57;
      11'd1366 : out_data_ref <= 8'h25;
      11'd1367 : out_data_ref <= 8'h29;
      11'd1368 : out_data_ref <= 8'h23;
      11'd1369 : out_data_ref <= 8'h8f;
      11'd1370 : out_data_ref <= 8'h92;
      11'd1371 : out_data_ref <= 8'hd3;
      11'd1372 : out_data_ref <= 8'hd8;
      11'd1373 : out_data_ref <= 8'hd2;
      11'd1374 : out_data_ref <= 8'hf3;
      11'd1375 : out_data_ref <= 8'hbc;
      11'd1376 : out_data_ref <= 8'hc5;
      11'd1377 : out_data_ref <= 8'h5f;
      11'd1378 : out_data_ref <= 8'h72;
      11'd1379 : out_data_ref <= 8'h77;
      11'd1380 : out_data_ref <= 8'h43;
      11'd1381 : out_data_ref <= 8'h00;
      11'd1382 : out_data_ref <= 8'h74;
      11'd1383 : out_data_ref <= 8'hd0;
      11'd1384 : out_data_ref <= 8'he7;
      11'd1385 : out_data_ref <= 8'h3d;
      11'd1386 : out_data_ref <= 8'h2d;
      11'd1387 : out_data_ref <= 8'h4a;
      11'd1388 : out_data_ref <= 8'hb9;
      11'd1389 : out_data_ref <= 8'h75;
      11'd1390 : out_data_ref <= 8'hb4;
      11'd1391 : out_data_ref <= 8'h7d;
      11'd1392 : out_data_ref <= 8'hd3;
      11'd1393 : out_data_ref <= 8'hd0;
      11'd1394 : out_data_ref <= 8'h77;
      11'd1395 : out_data_ref <= 8'ha9;
      11'd1396 : out_data_ref <= 8'hf4;
      11'd1397 : out_data_ref <= 8'ha8;
      11'd1398 : out_data_ref <= 8'h6b;
      11'd1399 : out_data_ref <= 8'h88;
      11'd1400 : out_data_ref <= 8'hdb;
      11'd1401 : out_data_ref <= 8'h44;
      11'd1402 : out_data_ref <= 8'h16;
      11'd1403 : out_data_ref <= 8'h69;
      11'd1404 : out_data_ref <= 8'h68;
      11'd1405 : out_data_ref <= 8'hee;
      11'd1406 : out_data_ref <= 8'h3d;
      11'd1407 : out_data_ref <= 8'hde;
      11'd1408 : out_data_ref <= 8'he1;
      11'd1409 : out_data_ref <= 8'h8b;
      11'd1410 : out_data_ref <= 8'h47;
      11'd1411 : out_data_ref <= 8'h2f;
      11'd1412 : out_data_ref <= 8'h93;
      11'd1413 : out_data_ref <= 8'hce;
      11'd1414 : out_data_ref <= 8'h05;
      11'd1415 : out_data_ref <= 8'he8;
      11'd1416 : out_data_ref <= 8'h19;
      11'd1417 : out_data_ref <= 8'h68;
      11'd1418 : out_data_ref <= 8'h72;
      11'd1419 : out_data_ref <= 8'hde;
      11'd1420 : out_data_ref <= 8'h78;
      11'd1421 : out_data_ref <= 8'h4c;
      11'd1422 : out_data_ref <= 8'hc9;
      11'd1423 : out_data_ref <= 8'h0a;
      11'd1424 : out_data_ref <= 8'hdc;
      11'd1425 : out_data_ref <= 8'h89;
      11'd1426 : out_data_ref <= 8'h00;
      11'd1427 : out_data_ref <= 8'h0d;
      11'd1428 : out_data_ref <= 8'h6c;
      11'd1429 : out_data_ref <= 8'hb9;
      11'd1430 : out_data_ref <= 8'h72;
      11'd1431 : out_data_ref <= 8'h1a;
      11'd1432 : out_data_ref <= 8'hc9;
      11'd1433 : out_data_ref <= 8'hf1;
      11'd1434 : out_data_ref <= 8'h36;
      11'd1435 : out_data_ref <= 8'h34;
      11'd1436 : out_data_ref <= 8'heb;
      11'd1437 : out_data_ref <= 8'he9;
      11'd1438 : out_data_ref <= 8'h8a;
      11'd1439 : out_data_ref <= 8'ha2;
      11'd1440 : out_data_ref <= 8'ha6;
      11'd1441 : out_data_ref <= 8'hdd;
      11'd1442 : out_data_ref <= 8'hee;
      11'd1443 : out_data_ref <= 8'h25;
      11'd1444 : out_data_ref <= 8'h39;
      11'd1445 : out_data_ref <= 8'hb5;
      11'd1446 : out_data_ref <= 8'h7f;
      11'd1447 : out_data_ref <= 8'hce;
      11'd1448 : out_data_ref <= 8'h84;
      11'd1449 : out_data_ref <= 8'hfc;
      11'd1450 : out_data_ref <= 8'h22;
      11'd1451 : out_data_ref <= 8'h08;
      11'd1452 : out_data_ref <= 8'h36;
      11'd1453 : out_data_ref <= 8'h5c;
      11'd1454 : out_data_ref <= 8'he2;
      11'd1455 : out_data_ref <= 8'h87;
      11'd1456 : out_data_ref <= 8'h2b;
      11'd1457 : out_data_ref <= 8'h35;
      11'd1458 : out_data_ref <= 8'hc2;
      11'd1459 : out_data_ref <= 8'h54;
      11'd1460 : out_data_ref <= 8'hf4;
      11'd1461 : out_data_ref <= 8'h8b;
      11'd1462 : out_data_ref <= 8'h4d;
      11'd1463 : out_data_ref <= 8'h9a;
      11'd1464 : out_data_ref <= 8'h32;
      11'd1465 : out_data_ref <= 8'h3f;
      11'd1466 : out_data_ref <= 8'h3f;
      11'd1467 : out_data_ref <= 8'h08;
      11'd1468 : out_data_ref <= 8'h6e;
      11'd1469 : out_data_ref <= 8'h20;
      11'd1470 : out_data_ref <= 8'hd9;
      11'd1471 : out_data_ref <= 8'ha2;
      11'd1472 : out_data_ref <= 8'hfc;
      11'd1473 : out_data_ref <= 8'he7;
      11'd1474 : out_data_ref <= 8'he5;
      11'd1475 : out_data_ref <= 8'hbe;
      11'd1476 : out_data_ref <= 8'hac;
      11'd1477 : out_data_ref <= 8'h80;
      11'd1478 : out_data_ref <= 8'h35;
      11'd1479 : out_data_ref <= 8'h32;
      11'd1480 : out_data_ref <= 8'hd9;
      11'd1481 : out_data_ref <= 8'h1e;
      11'd1482 : out_data_ref <= 8'hac;
      11'd1483 : out_data_ref <= 8'he6;
      11'd1484 : out_data_ref <= 8'h35;
      11'd1485 : out_data_ref <= 8'he8;
      11'd1486 : out_data_ref <= 8'h90;
      11'd1487 : out_data_ref <= 8'hbf;
      11'd1488 : out_data_ref <= 8'ha1;
      11'd1489 : out_data_ref <= 8'h14;
      11'd1490 : out_data_ref <= 8'h90;
      11'd1491 : out_data_ref <= 8'h77;
      11'd1492 : out_data_ref <= 8'h93;
      11'd1493 : out_data_ref <= 8'h99;
      11'd1494 : out_data_ref <= 8'hc0;
      11'd1495 : out_data_ref <= 8'h47;
      11'd1496 : out_data_ref <= 8'h6d;
      11'd1497 : out_data_ref <= 8'hdb;
      11'd1498 : out_data_ref <= 8'h0a;
      11'd1499 : out_data_ref <= 8'h87;
      11'd1500 : out_data_ref <= 8'hea;
      11'd1501 : out_data_ref <= 8'h54;
      11'd1502 : out_data_ref <= 8'h57;
      11'd1503 : out_data_ref <= 8'h55;
      11'd1504 : out_data_ref <= 8'hb0;
      11'd1505 : out_data_ref <= 8'h51;
      11'd1506 : out_data_ref <= 8'h43;
      11'd1507 : out_data_ref <= 8'hfb;
      11'd1508 : out_data_ref <= 8'h2e;
      11'd1509 : out_data_ref <= 8'ha1;
      11'd1510 : out_data_ref <= 8'h02;
      11'd1511 : out_data_ref <= 8'hfd;
      11'd1512 : out_data_ref <= 8'hf5;
      11'd1513 : out_data_ref <= 8'ha6;
      11'd1514 : out_data_ref <= 8'h54;
      11'd1515 : out_data_ref <= 8'h16;
      11'd1516 : out_data_ref <= 8'hfd;
      11'd1517 : out_data_ref <= 8'hae;
      11'd1518 : out_data_ref <= 8'h05;
      11'd1519 : out_data_ref <= 8'h65;
      11'd1520 : out_data_ref <= 8'h13;
      11'd1521 : out_data_ref <= 8'h37;
      11'd1522 : out_data_ref <= 8'hd6;
      11'd1523 : out_data_ref <= 8'hb6;
      11'd1524 : out_data_ref <= 8'h10;
      11'd1525 : out_data_ref <= 8'hcc;
      11'd1526 : out_data_ref <= 8'h85;
      11'd1527 : out_data_ref <= 8'h2b;
      11'd1528 : out_data_ref <= 8'h97;
      11'd1529 : out_data_ref <= 8'hc1;
      11'd1530 : out_data_ref <= 8'h82;
      11'd1531 : out_data_ref <= 8'h1f;
      11'd1532 : out_data_ref <= 8'h4c;
      11'd1533 : out_data_ref <= 8'hd3;
      11'd1534 : out_data_ref <= 8'hd6;
      11'd1535 : out_data_ref <= 8'heb;
      11'd1536 : out_data_ref <= 8'h95;
      11'd1537 : out_data_ref <= 8'h13;
      11'd1538 : out_data_ref <= 8'h2f;
      11'd1539 : out_data_ref <= 8'hb9;
      11'd1540 : out_data_ref <= 8'h4d;
      11'd1541 : out_data_ref <= 8'h62;
      11'd1542 : out_data_ref <= 8'h85;
      11'd1543 : out_data_ref <= 8'hd8;
      11'd1544 : out_data_ref <= 8'ha2;
      11'd1545 : out_data_ref <= 8'h39;
      11'd1546 : out_data_ref <= 8'h76;
      11'd1547 : out_data_ref <= 8'h87;
      11'd1548 : out_data_ref <= 8'hb0;
      11'd1549 : out_data_ref <= 8'h22;
      11'd1550 : out_data_ref <= 8'h0c;
      11'd1551 : out_data_ref <= 8'hc2;
      11'd1552 : out_data_ref <= 8'h55;
      11'd1553 : out_data_ref <= 8'ha8;
      11'd1554 : out_data_ref <= 8'h18;
      11'd1555 : out_data_ref <= 8'h06;
      11'd1556 : out_data_ref <= 8'hfa;
      11'd1557 : out_data_ref <= 8'he9;
      11'd1558 : out_data_ref <= 8'hd6;
      11'd1559 : out_data_ref <= 8'hee;
      11'd1560 : out_data_ref <= 8'hd8;
      11'd1561 : out_data_ref <= 8'h9c;
      11'd1562 : out_data_ref <= 8'h9f;
      11'd1563 : out_data_ref <= 8'haa;
      11'd1564 : out_data_ref <= 8'h1e;
      11'd1565 : out_data_ref <= 8'h42;
      11'd1566 : out_data_ref <= 8'ha9;
      11'd1567 : out_data_ref <= 8'ha5;
      11'd1568 : out_data_ref <= 8'h13;
      11'd1569 : out_data_ref <= 8'h3a;
      11'd1570 : out_data_ref <= 8'h4b;
      11'd1571 : out_data_ref <= 8'hd5;
      11'd1572 : out_data_ref <= 8'hf3;
      11'd1573 : out_data_ref <= 8'h21;
      11'd1574 : out_data_ref <= 8'hb9;
      11'd1575 : out_data_ref <= 8'h52;
      11'd1576 : out_data_ref <= 8'h3e;
      11'd1577 : out_data_ref <= 8'h82;
      11'd1578 : out_data_ref <= 8'h7a;
      11'd1579 : out_data_ref <= 8'h69;
      11'd1580 : out_data_ref <= 8'h63;
      11'd1581 : out_data_ref <= 8'h7b;
      11'd1582 : out_data_ref <= 8'h42;
      11'd1583 : out_data_ref <= 8'h89;
      11'd1584 : out_data_ref <= 8'h36;
      11'd1585 : out_data_ref <= 8'h7e;
      11'd1586 : out_data_ref <= 8'h91;
      11'd1587 : out_data_ref <= 8'h26;
      11'd1588 : out_data_ref <= 8'he8;
      11'd1589 : out_data_ref <= 8'h63;
      11'd1590 : out_data_ref <= 8'h29;
      11'd1591 : out_data_ref <= 8'hd4;
      11'd1592 : out_data_ref <= 8'h26;
      11'd1593 : out_data_ref <= 8'h69;
      11'd1594 : out_data_ref <= 8'h71;
      11'd1595 : out_data_ref <= 8'haa;
      11'd1596 : out_data_ref <= 8'he2;
      11'd1597 : out_data_ref <= 8'h86;
      11'd1598 : out_data_ref <= 8'h50;
      11'd1599 : out_data_ref <= 8'h68;
      11'd1600 : out_data_ref <= 8'h42;
      11'd1601 : out_data_ref <= 8'h4a;
      11'd1602 : out_data_ref <= 8'hb2;
      11'd1603 : out_data_ref <= 8'h06;
      11'd1604 : out_data_ref <= 8'ha0;
      11'd1605 : out_data_ref <= 8'h56;
      11'd1606 : out_data_ref <= 8'h5e;
      11'd1607 : out_data_ref <= 8'h48;
      11'd1608 : out_data_ref <= 8'h21;
      11'd1609 : out_data_ref <= 8'h88;
      11'd1610 : out_data_ref <= 8'h22;
      11'd1611 : out_data_ref <= 8'h89;
      11'd1612 : out_data_ref <= 8'h9b;
      11'd1613 : out_data_ref <= 8'ha2;
      11'd1614 : out_data_ref <= 8'hed;
      11'd1615 : out_data_ref <= 8'he6;
      11'd1616 : out_data_ref <= 8'he5;
      11'd1617 : out_data_ref <= 8'hb5;
      11'd1618 : out_data_ref <= 8'h7c;
      11'd1619 : out_data_ref <= 8'h9d;
      11'd1620 : out_data_ref <= 8'h8b;
      11'd1621 : out_data_ref <= 8'h4a;
      11'd1622 : out_data_ref <= 8'h00;
      default  : out_data_ref <= 8'h0;
    endcase
  end

endmodule
