module mod7177Svec35 (
    input       [34:0] z_in,
    output      [11:0] p0,
    output reg  [12:0] p1,
    output reg  [11:0] p2,
    output reg  [12:0] p3,
    output reg  [11:0] n0,
    output reg  [12:0] n1
) ;

    assign p0 = z_in[11:0];

    always @ (*) begin
        case({ z_in[26], z_in[24], z_in[18], z_in[15], z_in[12] })
            5'h00: p1 = 13'd0;
            5'h01: p1 = 13'd4096;
            5'h02: p1 = 13'd4060;
            5'h03: p1 = 13'd979;
            5'h04: p1 = 13'd3772;
            5'h05: p1 = 13'd691;
            5'h06: p1 = 13'd655;
            5'h07: p1 = 13'd4751;
            5'h08: p1 = 13'd4567;
            5'h09: p1 = 13'd1486;
            5'h0a: p1 = 13'd1450;
            5'h0b: p1 = 13'd5546;
            5'h0c: p1 = 13'd1162;
            5'h0d: p1 = 13'd5258;
            5'h0e: p1 = 13'd5222;
            5'h0f: p1 = 13'd2141;
            5'h10: p1 = 13'd3914;
            5'h11: p1 = 13'd833;
            5'h12: p1 = 13'd797;
            5'h13: p1 = 13'd4893;
            5'h14: p1 = 13'd509;
            5'h15: p1 = 13'd4605;
            5'h16: p1 = 13'd4569;
            5'h17: p1 = 13'd1488;
            5'h18: p1 = 13'd1304;
            5'h19: p1 = 13'd5400;
            5'h1a: p1 = 13'd5364;
            5'h1b: p1 = 13'd2283;
            5'h1c: p1 = 13'd5076;
            5'h1d: p1 = 13'd1995;
            5'h1e: p1 = 13'd1959;
            5'h1f: p1 = 13'd6055;
        endcase
    end

    always @ (*) begin
        case({ z_in[27], z_in[20], z_in[19], z_in[16], z_in[13] })
            5'h00: p2 = 12'd0;
            5'h01: p2 = 12'd1015;
            5'h02: p2 = 12'd943;
            5'h03: p2 = 12'd1958;
            5'h04: p2 = 12'd367;
            5'h05: p2 = 12'd1382;
            5'h06: p2 = 12'd1310;
            5'h07: p2 = 12'd2325;
            5'h08: p2 = 12'd734;
            5'h09: p2 = 12'd1749;
            5'h0a: p2 = 12'd1677;
            5'h0b: p2 = 12'd2692;
            5'h0c: p2 = 12'd1101;
            5'h0d: p2 = 12'd2116;
            5'h0e: p2 = 12'd2044;
            5'h0f: p2 = 12'd3059;
            5'h10: p2 = 12'd651;
            5'h11: p2 = 12'd1666;
            5'h12: p2 = 12'd1594;
            5'h13: p2 = 12'd2609;
            5'h14: p2 = 12'd1018;
            5'h15: p2 = 12'd2033;
            5'h16: p2 = 12'd1961;
            5'h17: p2 = 12'd2976;
            5'h18: p2 = 12'd1385;
            5'h19: p2 = 12'd2400;
            5'h1a: p2 = 12'd2328;
            5'h1b: p2 = 12'd3343;
            5'h1c: p2 = 12'd1752;
            5'h1d: p2 = 12'd2767;
            5'h1e: p2 = 12'd2695;
            5'h1f: p2 = 12'd3710;
        endcase
    end

    always @ (*) begin
        case({ z_in[34], z_in[31], z_in[30], z_in[29], z_in[22] })
            5'h00: p3 = 13'd0;
            5'h01: p3 = 13'd2936;
            5'h02: p3 = 13'd2604;
            5'h03: p3 = 13'd5540;
            5'h04: p3 = 13'd5208;
            5'h05: p3 = 13'd967;
            5'h06: p3 = 13'd635;
            5'h07: p3 = 13'd3571;
            5'h08: p3 = 13'd3239;
            5'h09: p3 = 13'd6175;
            5'h0a: p3 = 13'd5843;
            5'h0b: p3 = 13'd1602;
            5'h0c: p3 = 13'd1270;
            5'h0d: p3 = 13'd4206;
            5'h0e: p3 = 13'd3874;
            5'h0f: p3 = 13'd6810;
            5'h10: p3 = 13'd2796;
            5'h11: p3 = 13'd5732;
            5'h12: p3 = 13'd5400;
            5'h13: p3 = 13'd1159;
            5'h14: p3 = 13'd827;
            5'h15: p3 = 13'd3763;
            5'h16: p3 = 13'd3431;
            5'h17: p3 = 13'd6367;
            5'h18: p3 = 13'd6035;
            5'h19: p3 = 13'd1794;
            5'h1a: p3 = 13'd1462;
            5'h1b: p3 = 13'd4398;
            5'h1c: p3 = 13'd4066;
            5'h1d: p3 = 13'd7002;
            5'h1e: p3 = 13'd6670;
            5'h1f: p3 = 13'd2429;
        endcase
    end

    always @ (*) begin
        case({ z_in[33], z_in[32], z_in[23] })
            3'h0: n0 = 12'd0;
            3'h1: n0 = 12'd1305;
            3'h2: n0 = 12'd699;
            3'h3: n0 = 12'd2004;
            3'h4: n0 = 12'd1398;
            3'h5: n0 = 12'd2703;
            3'h6: n0 = 12'd2097;
            3'h7: n0 = 12'd3402;
        endcase
    end

    always @ (*) begin
        case({ z_in[28], z_in[25], z_in[21], z_in[17], z_in[14] })
            5'h00: n1 = 13'd0;
            5'h01: n1 = 13'd5147;
            5'h02: n1 = 13'd5291;
            5'h03: n1 = 13'd3261;
            5'h04: n1 = 13'd5709;
            5'h05: n1 = 13'd3679;
            5'h06: n1 = 13'd3823;
            5'h07: n1 = 13'd1793;
            5'h08: n1 = 13'd5220;
            5'h09: n1 = 13'd3190;
            5'h0a: n1 = 13'd3334;
            5'h0b: n1 = 13'd1304;
            5'h0c: n1 = 13'd3752;
            5'h0d: n1 = 13'd1722;
            5'h0e: n1 = 13'd1866;
            5'h0f: n1 = 13'd7013;
            5'h10: n1 = 13'd5875;
            5'h11: n1 = 13'd3845;
            5'h12: n1 = 13'd3989;
            5'h13: n1 = 13'd1959;
            5'h14: n1 = 13'd4407;
            5'h15: n1 = 13'd2377;
            5'h16: n1 = 13'd2521;
            5'h17: n1 = 13'd491;
            5'h18: n1 = 13'd3918;
            5'h19: n1 = 13'd1888;
            5'h1a: n1 = 13'd2032;
            5'h1b: n1 = 13'd2;
            5'h1c: n1 = 13'd2450;
            5'h1d: n1 = 13'd420;
            5'h1e: n1 = 13'd564;
            5'h1f: n1 = 13'd5711;
        endcase
    end

endmodule
