module ntt4096_163841 ( clk, rst, start, input_fg, addr, din, dout, valid );

  localparam Q0 = 163841;

  // STATE
  localparam ST_IDLE   = 0;
  localparam ST_NTT    = 1;
  localparam ST_PMUL   = 2;
  localparam ST_RELOAD = 3;
  localparam ST_INTT   = 4;
  localparam ST_CRT    = 5;  // not applied for single prime scheme
  localparam ST_REDUCE = 6;
  localparam ST_FINISH = 7;

  input                      clk;
  input                      rst;
  input                      start;
  input                      input_fg;
  input             [12 : 0] addr;
  input signed      [17 : 0] din;
  output reg signed [17 : 0] dout;
  output reg                 valid;

  // BRAM
  reg            wr_en   [0 : 1];
  reg   [12 : 0] wr_addr [0 : 1];
  reg   [12 : 0] rd_addr [0 : 1];
  reg   [17 : 0] wr_din  [0 : 1];
  wire  [17 : 0] rd_dout [0 : 1];
  wire  [17 : 0] wr_dout [0 : 1];

  // addr_gen
  wire         bank_index_rd [0 : 1];
  wire         bank_index_wr [0 : 1];
  wire [11: 0] data_index_rd [0 : 1];
  wire [11: 0] data_index_wr [0 : 1];
  reg  bank_index_wr_0_shift_1, bank_index_wr_0_shift_2;
  reg  fg_shift_1, fg_shift_2, fg_shift_3;

  // w_addr_gen
  reg  [11 : 0] stage_bit;
  wire [11 : 0] w_addr;

  // bfu
  reg                  ntt_state; 
  reg  signed [17: 0] in_a  ;
  reg  signed [17: 0] in_b  ;
  reg  signed [17: 0] in_w  ;
  wire signed [35: 0] bw    ;
  wire signed [17: 0] out_a ;
  wire signed [17: 0] out_b ;

  // state, stage, counter
  reg  [2 : 0] state, next_state;
  reg  [4 : 0] stage, stage_wr;
  wire [4 : 0] stage_rdM, stage_wrM;
  reg  [13 : 0] ctr;
  reg  [13 : 0] ctr_shift_7, ctr_shift_8, ctr_shift_9, ctr_shift_1, ctr_shift_2;
  reg          ctr_MSB_masked;
  reg          poly_select;
  reg          ctr_msb_shift_1;
  wire         ctr_half_end, ctr_full_end, ctr_shift_7_end, stage_rd_end, stage_rd_2, stage_wr_end, ntt_end, point_proc_end, reduce_end;

  // w_array
  reg         [12: 0] w_addr_in;
  wire signed [17: 0] w_dout ;

  // misc
  reg          bank_index_rd_shift_1, bank_index_rd_shift_2;
  reg [12: 0] wr_ctr [0 : 1];
  reg [17: 0] din_shift_1, din_shift_2, din_shift_3;
  reg [12: 0] w_addr_in_shift_1;

  // BRAM instances
  bram_18_13_P bank_0
  (clk, wr_en[0], wr_addr[0], rd_addr[0], wr_din[0], wr_dout[0], rd_dout[0]);
  bram_18_13_P bank_1
  (clk, wr_en[1], wr_addr[1], rd_addr[1], wr_din[1], wr_dout[1], rd_dout[1]);

  // Read/Write Address Generator
  addr_gen addr_rd_0 (clk, stage_rdM, {ctr_MSB_masked, ctr[11:0]}, bank_index_rd[0], data_index_rd[0]);
  addr_gen addr_rd_1 (clk, stage_rdM, {1'b1, ctr[11:0]}, bank_index_rd[1], data_index_rd[1]);
  addr_gen addr_wr_0 (clk, stage_wrM, {wr_ctr[0]}, bank_index_wr[0], data_index_wr[0]);
  addr_gen addr_wr_1 (clk, stage_wrM, {wr_ctr[1]}, bank_index_wr[1], data_index_wr[1]);

  // Omega Address Generator
  w_addr_gen w_addr_gen_0 (clk, stage_bit, ctr[11:0], w_addr);

  // Butterfly Unit  , each with a corresponding omega array
  bfu_163841 bfu_inst (clk, ntt_state, in_a, in_b, in_w, bw, out_a, out_b);
  w_163841 rom_w_inst (clk, w_addr_in_shift_1, w_dout);

  assign ctr_half_end         = (ctr[11:0] == 4095) ? 1 : 0;
  assign ctr_full_end         = (ctr[12:0] == 8191) ? 1 : 0;
  assign stage_rd_end         = (stage == 13) ? 1 : 0;
  assign stage_rd_2           = (stage == 2) ? 1 : 0;
  assign ntt_end         = (stage_rd_end && ctr[11 : 0] == 10) ? 1 : 0;
  assign crt_end         = (stage_rd_2 && ctr[11 : 0] == 10) ? 1 : 0;
  assign point_proc_end   = (ctr == 8202) ? 1 : 0;
  assign reload_end      = (stage != 0 && ctr[11:0] == 4) ? 1 : 0;
  assign reduce_end      = (ctr == 8196);

  // crt
  // fg_shift
  always @ ( posedge clk ) begin
    fg_shift_1 <= input_fg;
    fg_shift_2 <= fg_shift_1;
    fg_shift_3 <= fg_shift_2;
  end
  // dout
  always @ ( posedge clk ) begin
    if (state == ST_FINISH) begin
      if (bank_index_wr_0_shift_2) begin
        dout <= wr_dout[1][17:0];
      end else begin
        dout <= wr_dout[0][17:0];
      end
    end else begin
      dout <= 'sd0;
    end
  end

  // bank_index_wr_0_shift_1
  always @ ( posedge clk ) begin
    bank_index_wr_0_shift_1 <= bank_index_wr[0];
    bank_index_wr_0_shift_2 <= bank_index_wr_0_shift_1;
  end

  // poly_select
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        poly_select <= ~poly_select;
      end else begin
        poly_select <= poly_select;
      end    
    end else if (state == ST_RELOAD) begin
      poly_select <= 1;
    end else begin
      poly_select <= 0;
    end
  end

  // w_addr_in_shift_1
  always @ ( posedge clk ) begin
    w_addr_in_shift_1 <= w_addr_in;
  end

  // din_shift
  always @ ( posedge clk ) begin
    din_shift_1 <= din;
    din_shift_2 <= din_shift_1;
    din_shift_3 <= din_shift_2;
  end

  // rd_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_rd[0]) begin
        rd_addr[0][11:0] <= data_index_rd[1];
        rd_addr[1][11:0] <= data_index_rd[0];
      end else begin
        rd_addr[0][11:0] <= data_index_rd[0];
        rd_addr[1][11:0] <= data_index_rd[1];
      end
    end else begin
      rd_addr[0][11:0] <= data_index_rd[0];
      rd_addr[1][11:0] <= data_index_rd[0];
    end

    if (state == ST_NTT)  begin
      rd_addr[0][12] <= poly_select;
      rd_addr[1][12] <= poly_select;
    end else if (state == ST_PMUL) begin
      rd_addr[0][12] <=  bank_index_rd[0];
      rd_addr[1][12] <= ~bank_index_rd[0];
    end else if (state == ST_RELOAD) begin
      rd_addr[0][12] <= 0;
      rd_addr[1][12] <= 0;
    end else begin
      rd_addr[0][12] <= 1;
      rd_addr[1][12] <= 1;
    end
  end

  // wr_en
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 1;
      end
    end else if (state == ST_IDLE) begin
      if (fg_shift_3 ^ bank_index_wr[0]) begin
        wr_en[0] <= 0;
        wr_en[1] <= 1;
      end else begin
        wr_en[0] <= 1;
        wr_en[1] <= 0;
      end
    end else if (state == ST_PMUL) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_REDUCE) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <= ~bank_index_wr[0];
        wr_en[1] <=  bank_index_wr[0];
      end
    end else if (state == ST_CRT) begin
      if (stage == 0 && ctr < 11) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else if (state == ST_RELOAD) begin
      if (stage == 0 && ctr < 4) begin
        wr_en[0] <= 0;
        wr_en[1] <= 0;
      end else begin
        wr_en[0] <=  bank_index_wr[0];
        wr_en[1] <= ~bank_index_wr[0];
      end
    end else begin
      wr_en[0] <= 0;
      wr_en[1] <= 0;
    end
  end

  // wr_addr
  always @(posedge clk ) begin
    if ( state == ST_NTT || state == ST_INTT ) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_addr[0][11:0] <= data_index_wr[1];
        wr_addr[1][11:0] <= data_index_wr[0];
      end else begin
        wr_addr[0][11:0] <= data_index_wr[0];
        wr_addr[1][11:0] <= data_index_wr[1];
      end
    end else begin
      wr_addr[0][11:0] <= data_index_wr[0];
      wr_addr[1][11:0] <= data_index_wr[0];
    end  

    if (state == ST_IDLE) begin
      wr_addr[0][12] <= fg_shift_3;
      wr_addr[1][12] <= fg_shift_3;
    end else if(state == ST_NTT || state == ST_INTT) begin
      wr_addr[0][12] <= poly_select;
      wr_addr[1][12] <= poly_select;
    end else if (state == ST_PMUL || state == ST_REDUCE || state == ST_FINISH) begin
      wr_addr[0][12] <= 0;
      wr_addr[1][12] <= 0;
    end else begin
      wr_addr[0][12] <= 1;
      wr_addr[1][12] <= 1;
    end     
  end

  // wr_din
  always @ ( posedge clk ) begin
    if (state == ST_IDLE) begin
      wr_din[0][17:0] <= { din_shift_3 };
      wr_din[1][17:0] <= { din_shift_3 };
    end else if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_wr[0]) begin
        wr_din[0][17:0] <= out_b;
        wr_din[1][17:0] <= out_a;
      end else begin
        wr_din[0][17:0] <= out_a;
        wr_din[1][17:0] <= out_b;
      end
    end else if (state == ST_RELOAD) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end
    end else if (state == ST_REDUCE) begin
      if (bank_index_rd_shift_2) begin
        wr_din[0][17:0] <= rd_dout[0][17:0];
        wr_din[1][17:0] <= rd_dout[0][17:0];
      end else begin
        wr_din[0][17:0] <= rd_dout[1][17:0];
        wr_din[1][17:0] <= rd_dout[1][17:0];
      end
    end else begin
      wr_din[0][17:0] <= out_a;
      wr_din[1][17:0] <= out_a;
    end
  end

  // bank_index_rd_shift
  always @ ( posedge clk ) begin
    bank_index_rd_shift_1 <= bank_index_rd[0];
    bank_index_rd_shift_2 <= bank_index_rd_shift_1;
  end

  // ntt_state
  always @ ( posedge clk ) begin
    if (state == ST_INTT) begin
      ntt_state <= 1;
    end else begin
      ntt_state <= 0;
    end
  end

  // in_a, in_b
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else if (state == ST_CRT) begin
      if (bank_index_rd_shift_2) begin
        in_b <= $signed(rd_dout[0]);
      end else begin
        in_b <= $signed(rd_dout[1]);
      end
    end else begin // ST_PMUL
      in_b <= $signed(rd_dout[1]);
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (poly_select ^ bank_index_rd_shift_2) begin
        in_a <= $signed(rd_dout[1]);
      end else begin
        in_a <= $signed(rd_dout[0]);
      end
    end else begin // ST_PMUL, ST_CRT
      in_a <= 'sd0;
    end
  end

  // w_addr_in, in_w
  always @ ( posedge clk ) begin
    if (state == ST_NTT) begin
      w_addr_in <= {1'b0, w_addr};
    end else begin
      w_addr_in <= 8192 - w_addr;
    end

    if (state == ST_PMUL) begin
        in_w <= rd_dout[0];
    end else begin
      in_w <= w_dout;
    end
  end

  // wr_ctr
  always @ ( posedge clk ) begin
    if (state == ST_IDLE || state == ST_FINISH) begin
      wr_ctr[0] <= addr[12:0];
    end else if (state == ST_RELOAD || state == ST_REDUCE) begin
      wr_ctr[0] <= {ctr_shift_1[0], ctr_shift_1[1], ctr_shift_1[2], ctr_shift_1[3], ctr_shift_1[4], ctr_shift_1[5], ctr_shift_1[6], ctr_shift_1[7], ctr_shift_1[8], ctr_shift_1[9], ctr_shift_1[10], ctr_shift_1[11], ctr_shift_1[12]};
    end else if (state == ST_NTT || state == ST_INTT) begin
      wr_ctr[0] <= {1'b0, ctr_shift_7[11:0]};
    end else begin
      wr_ctr[0] <= ctr_shift_7[12:0];
    end

    wr_ctr[1] <= {1'b1, ctr_shift_7[11:0]};
  end

  // ctr_MSB_masked
  always @ (*) begin
    if (state == ST_NTT || state == ST_INTT) begin
      ctr_MSB_masked = 0;
    end else begin
      ctr_MSB_masked = ctr[12];
    end
  end

  // ctr, ctr_shifts
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_PMUL) begin
      if (point_proc_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_CRT) begin
      if (crt_end || ctr_full_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else if (state == ST_REDUCE) begin
      if (reduce_end) begin
        ctr <= 0;
      end else begin
        ctr <= ctr + 1;
      end
    end else begin
      ctr <= 0;
    end

    //change ctr_shift_7 <= ctr - 5;
    ctr_shift_7 <= ctr - 7;
    ctr_shift_8 <= ctr_shift_7;
    ctr_shift_9 <= ctr_shift_8;
    ctr_shift_1 <= ctr;
    ctr_shift_2 <= ctr_shift_1;
  end

  // stage, stage_wr
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage <= 0;
      end else if (ctr_half_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage <= 0;
      end else if (ctr_full_end) begin
        stage <= stage + 1;
      end else begin
        stage <= stage;
      end
    end else begin
      stage <= 0;
    end

    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[11:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_RELOAD) begin
      if (reload_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_7[12:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else if (state == ST_CRT) begin
      if (crt_end) begin
        stage_wr <= 0;
      end else if (ctr_shift_9[12:0] == 0 && stage != 0) begin
        stage_wr <= stage_wr + 1;
      end else begin
        stage_wr <= stage_wr;
      end
    end else begin
      stage_wr <= 0;
    end        
  end
  assign stage_rdM = (state == ST_NTT || state == ST_INTT) ? stage : 0;
  assign stage_wrM = (state == ST_NTT || state == ST_INTT) ? stage_wr : 0;

  // stage_bit
  always @ ( posedge clk ) begin
    if (state == ST_NTT || state == ST_INTT) begin
      if (ntt_end) begin
        stage_bit <= 0;
      end else if (ctr_half_end) begin
        stage_bit[0] <= 1'b1;
        stage_bit[11 : 1] <= stage_bit[10 : 0];
      end else begin
        stage_bit <= stage_bit;
      end
    end else begin
      stage_bit <= 'b0;
    end
  end

  // valid
  always @ (*) begin
      if (state == ST_FINISH) begin
          valid = 1;
      end else begin
          valid = 0;
      end
  end

  // state
  always @ ( posedge clk ) begin
    if(rst) begin
            state <= 0;
        end else begin
            state <= next_state;
        end
  end

  always @(*) begin
    case(state)
    ST_IDLE: begin
      if(start)
        next_state = ST_NTT;
      else
        next_state = ST_IDLE;
    end
    ST_NTT: begin
      if(ntt_end && poly_select == 1)
        next_state = ST_PMUL;
      else
        next_state = ST_NTT;
    end
    ST_PMUL: begin
      if (point_proc_end)
        next_state = ST_RELOAD;
      else
        next_state = ST_PMUL;
    end
    ST_RELOAD: begin
      if (reload_end) begin
        next_state = ST_INTT;
      end else begin
        next_state = ST_RELOAD;
      end
    end
    ST_INTT: begin
      if(ntt_end)
        next_state = ST_REDUCE;
      else
        next_state = ST_INTT;
      end
    ST_REDUCE: begin
      if(reduce_end)
        next_state = ST_FINISH;
      else
        next_state = ST_REDUCE;
    end
    ST_FINISH: begin
      if(!start)
        next_state = ST_FINISH;
      else
        next_state = ST_IDLE;
    end
    default: next_state = ST_IDLE;
    endcase
  end

endmodule

module w_addr_gen ( clk, stage_bit, ctr, w_addr );

  input              clk;
  input      [11: 0] stage_bit;
  input      [11: 0] ctr;
  output reg [11: 0] w_addr;

  wire [11: 0] w;

  assign w[ 0] = (stage_bit[ 0]) ? ctr[ 0] : 0;
  assign w[ 1] = (stage_bit[ 1]) ? ctr[ 1] : 0;
  assign w[ 2] = (stage_bit[ 2]) ? ctr[ 2] : 0;
  assign w[ 3] = (stage_bit[ 3]) ? ctr[ 3] : 0;
  assign w[ 4] = (stage_bit[ 4]) ? ctr[ 4] : 0;
  assign w[ 5] = (stage_bit[ 5]) ? ctr[ 5] : 0;
  assign w[ 6] = (stage_bit[ 6]) ? ctr[ 6] : 0;
  assign w[ 7] = (stage_bit[ 7]) ? ctr[ 7] : 0;
  assign w[ 8] = (stage_bit[ 8]) ? ctr[ 8] : 0;
  assign w[ 9] = (stage_bit[ 9]) ? ctr[ 9] : 0;
  assign w[10] = (stage_bit[10]) ? ctr[10] : 0;
  assign w[11] = (stage_bit[11]) ? ctr[11] : 0;

  always @ ( posedge clk ) begin
    w_addr <= {w[0], w[1], w[2], w[3], w[4], w[5], w[6], w[7], w[8], w[9], w[10], w[11]};
  end

endmodule

module addr_gen ( clk, stage, ctr, bank_index, data_index );

  input              clk;
  input      [3 : 0] stage;
  input      [12: 0] ctr;
  output reg         bank_index;
  output reg [11: 0] data_index;

  wire       [12: 0] bs_out;

  barrel_shifter bs ( clk, ctr, stage, bs_out );

    always @( posedge clk ) begin
        bank_index <= ^bs_out;
    end

    always @( posedge clk ) begin
        data_index <= bs_out[12:1];
    end

endmodule

module barrel_shifter ( clk, in, shift, out );

  input              clk;
  input      [12: 0] in;
  input      [3 : 0] shift;
  output reg [12: 0] out;

  reg        [12: 0] in_s [0:4];

  always @ (*) begin
    in_s[0] = in;
  end

  always @ (*) begin
    if(shift[0]) begin
      in_s[1] = { in_s[0][0], in_s[0][12:1] };
    end else begin
      in_s[1] = in_s[0];
    end
  end

  always @ (*) begin
    if(shift[1]) begin
      in_s[2] = { in_s[1][1:0], in_s[1][12:2] };
    end else begin
      in_s[2] = in_s[1];
    end
  end

  always @ (*) begin
    if(shift[2]) begin
      in_s[3] = { in_s[2][3:0], in_s[2][12:4] };
    end else begin
      in_s[3] = in_s[2];
    end
  end

  always @ (*) begin
    if(shift[3]) begin
      in_s[4] = { in_s[3][7:0], in_s[3][12:8] };
    end else begin
      in_s[4] = in_s[3];
    end
  end

  always @ ( posedge clk ) begin
    out <= in_s[4];
  end

endmodule

module bfu_163841 ( clk, state, in_a, in_b, w, bw, out_a, out_b );

  input                      clk;
  input                      state;
  input      signed [17 : 0] in_a;
  input      signed [17 : 0] in_b;
  input      signed [17 : 0] w;
  output reg signed [34 : 0] bw;
  output reg signed [17 : 0] out_a;
  output reg signed [17 : 0] out_b;

  wire signed       [17 : 0] mod_bw;
  reg signed        [18 : 0] a, b;
  reg signed        [17 : 0] in_a_s1, in_a_s2, in_a_s3, in_a_s4, in_a_s5;

  reg signed        [34 : 0] bwQ_0, bwQ_1, bwQ_2;
  wire signed       [18 : 0] a_add_q, a_sub_q, b_add_q, b_sub_q;

  modmul163841s mod163841s_inst ( clk, 1'b0, bw, mod_bw );

  assign a_add_q = a + 'sd163841;
  assign a_sub_q = a - 'sd163841;
  assign b_add_q = b + 'sd163841;
  assign b_sub_q = b - 'sd163841;

  always @(posedge clk ) begin
    in_a_s1 <= in_a;
    in_a_s2 <= in_a_s1;
    in_a_s3 <= in_a_s2;
    in_a_s4 <= in_a_s3;
    in_a_s5 <= in_a_s4;
  end

  always @ ( posedge clk ) begin
    bw <= in_b * w;
  end

  always @ ( posedge clk ) begin
    a <= in_a_s4 + mod_bw;
    b <= in_a_s4 - mod_bw;

    if (state == 0) begin
      if (a > 'sd81920) begin
        out_a <= a_sub_q;
      end else if (a < -'sd81920) begin
        out_a <= a_add_q;
      end else begin
        out_a <= a;
      end
    end else begin
      if (a[0] == 0) begin
        out_a <= a[18:1];
      end else if (a[18] == 0) begin // a > 0
        out_a <= a_sub_q[18:1];
      end else begin                 // a < 0
        out_a <= a_add_q[18:1];
      end
    end

    if (state == 0) begin
      if (b > 'sd81920) begin
        out_b <= b_sub_q;
      end else if (b < -'sd81920) begin
        out_b <= b_add_q;
      end else begin
        out_b <= b;
      end
    end else begin
      if (b[0] == 0) begin
        out_b <= b[18:1];
      end else if (b[18] == 0) begin // b > 0
        out_b <= b_sub_q[18:1];
      end else begin                 // b < 0
        out_b <= b_add_q[18:1];
      end
    end
  end

endmodule

module w_163841 ( clk, addr, dout );

  input                       clk;
  input             [12 : 0]  addr;
  output signed     [17 : 0]  dout;

  wire signed       [17 : 0]  dout_p;
  wire signed       [17 : 0]  dout_n;
  reg               [12 : 0]  addr_reg;

  (* rom_style = "block" *) reg signed [17:0] data [0:4095];

  assign dout_p = data[addr_reg[11:0]];
  assign dout_n = -dout_p;
  assign dout   = addr_reg[12] ? dout_n : dout_p;

  always @ ( posedge clk ) begin
    addr_reg <= addr;
  end

  initial begin
    data[   0] =  'sd1;
    data[   1] =  'sd25;
    data[   2] =  'sd625;
    data[   3] =  'sd15625;
    data[   4] =  'sd62943;
    data[   5] = -'sd64835;
    data[   6] =  'sd17535;
    data[   7] = -'sd53148;
    data[   8] = -'sd17972;
    data[   9] =  'sd42223;
    data[  10] =  'sd72529;
    data[  11] =  'sd10974;
    data[  12] = -'sd53332;
    data[  13] = -'sd22572;
    data[  14] = -'sd72777;
    data[  15] = -'sd17174;
    data[  16] =  'sd62173;
    data[  17] =  'sd79756;
    data[  18] =  'sd27808;
    data[  19] =  'sd39836;
    data[  20] =  'sd12854;
    data[  21] = -'sd6332;
    data[  22] =  'sd5541;
    data[  23] = -'sd25316;
    data[  24] =  'sd22464;
    data[  25] =  'sd70077;
    data[  26] = -'sd50326;
    data[  27] =  'sd52578;
    data[  28] =  'sd3722;
    data[  29] = -'sd70791;
    data[  30] =  'sd32476;
    data[  31] = -'sd7305;
    data[  32] = -'sd18784;
    data[  33] =  'sd21923;
    data[  34] =  'sd56552;
    data[  35] = -'sd60769;
    data[  36] = -'sd44656;
    data[  37] =  'sd30487;
    data[  38] = -'sd57030;
    data[  39] =  'sd48819;
    data[  40] =  'sd73588;
    data[  41] =  'sd37449;
    data[  42] = -'sd46821;
    data[  43] = -'sd23638;
    data[  44] =  'sd64414;
    data[  45] = -'sd28060;
    data[  46] = -'sd46136;
    data[  47] = -'sd6513;
    data[  48] =  'sd1016;
    data[  49] =  'sd25400;
    data[  50] = -'sd20364;
    data[  51] = -'sd17577;
    data[  52] =  'sd52098;
    data[  53] = -'sd8278;
    data[  54] = -'sd43109;
    data[  55] =  'sd69162;
    data[  56] = -'sd73201;
    data[  57] = -'sd27774;
    data[  58] = -'sd38986;
    data[  59] =  'sd8396;
    data[  60] =  'sd46059;
    data[  61] =  'sd4588;
    data[  62] = -'sd49141;
    data[  63] = -'sd81638;
    data[  64] = -'sd74858;
    data[  65] = -'sd69199;
    data[  66] =  'sd72276;
    data[  67] =  'sd4649;
    data[  68] = -'sd47616;
    data[  69] = -'sd43513;
    data[  70] =  'sd59062;
    data[  71] =  'sd1981;
    data[  72] =  'sd49525;
    data[  73] = -'sd72603;
    data[  74] = -'sd12824;
    data[  75] =  'sd7082;
    data[  76] =  'sd13209;
    data[  77] =  'sd2543;
    data[  78] =  'sd63575;
    data[  79] = -'sd49035;
    data[  80] = -'sd78988;
    data[  81] = -'sd8608;
    data[  82] = -'sd51359;
    data[  83] =  'sd26753;
    data[  84] =  'sd13461;
    data[  85] =  'sd8843;
    data[  86] =  'sd57234;
    data[  87] = -'sd43719;
    data[  88] =  'sd53912;
    data[  89] =  'sd37072;
    data[  90] = -'sd56246;
    data[  91] =  'sd68419;
    data[  92] =  'sd72065;
    data[  93] = -'sd626;
    data[  94] = -'sd15650;
    data[  95] = -'sd63568;
    data[  96] =  'sd49210;
    data[  97] = -'sd80478;
    data[  98] = -'sd45858;
    data[  99] =  'sd437;
    data[ 100] =  'sd10925;
    data[ 101] = -'sd54557;
    data[ 102] = -'sd53197;
    data[ 103] = -'sd19197;
    data[ 104] =  'sd11598;
    data[ 105] = -'sd37732;
    data[ 106] =  'sd39746;
    data[ 107] =  'sd10604;
    data[ 108] = -'sd62582;
    data[ 109] =  'sd73860;
    data[ 110] =  'sd44249;
    data[ 111] = -'sd40662;
    data[ 112] = -'sd33504;
    data[ 113] = -'sd18395;
    data[ 114] =  'sd31648;
    data[ 115] = -'sd28005;
    data[ 116] = -'sd44761;
    data[ 117] =  'sd27862;
    data[ 118] =  'sd41186;
    data[ 119] =  'sd46604;
    data[ 120] =  'sd18213;
    data[ 121] = -'sd36198;
    data[ 122] =  'sd78096;
    data[ 123] = -'sd13692;
    data[ 124] = -'sd14618;
    data[ 125] = -'sd37768;
    data[ 126] =  'sd38846;
    data[ 127] = -'sd11896;
    data[ 128] =  'sd30282;
    data[ 129] = -'sd62155;
    data[ 130] = -'sd79306;
    data[ 131] = -'sd16558;
    data[ 132] =  'sd77573;
    data[ 133] = -'sd26767;
    data[ 134] = -'sd13811;
    data[ 135] = -'sd17593;
    data[ 136] =  'sd51698;
    data[ 137] = -'sd18278;
    data[ 138] =  'sd34573;
    data[ 139] =  'sd45120;
    data[ 140] = -'sd18887;
    data[ 141] =  'sd19348;
    data[ 142] = -'sd7823;
    data[ 143] = -'sd31734;
    data[ 144] =  'sd25855;
    data[ 145] = -'sd8989;
    data[ 146] = -'sd60884;
    data[ 147] = -'sd47531;
    data[ 148] = -'sd41388;
    data[ 149] = -'sd51654;
    data[ 150] =  'sd19378;
    data[ 151] = -'sd7073;
    data[ 152] = -'sd12984;
    data[ 153] =  'sd3082;
    data[ 154] =  'sd77050;
    data[ 155] = -'sd39842;
    data[ 156] = -'sd13004;
    data[ 157] =  'sd2582;
    data[ 158] =  'sd64550;
    data[ 159] = -'sd24660;
    data[ 160] =  'sd38864;
    data[ 161] = -'sd11446;
    data[ 162] =  'sd41532;
    data[ 163] =  'sd55254;
    data[ 164] =  'sd70622;
    data[ 165] = -'sd36701;
    data[ 166] =  'sd65521;
    data[ 167] = -'sd385;
    data[ 168] = -'sd9625;
    data[ 169] = -'sd76784;
    data[ 170] =  'sd46492;
    data[ 171] =  'sd15413;
    data[ 172] =  'sd57643;
    data[ 173] = -'sd33494;
    data[ 174] = -'sd18145;
    data[ 175] =  'sd37898;
    data[ 176] = -'sd35596;
    data[ 177] = -'sd70695;
    data[ 178] =  'sd34876;
    data[ 179] =  'sd52695;
    data[ 180] =  'sd6647;
    data[ 181] =  'sd2334;
    data[ 182] =  'sd58350;
    data[ 183] = -'sd15819;
    data[ 184] = -'sd67793;
    data[ 185] = -'sd56415;
    data[ 186] =  'sd64194;
    data[ 187] = -'sd33560;
    data[ 188] = -'sd19795;
    data[ 189] = -'sd3352;
    data[ 190] =  'sd80041;
    data[ 191] =  'sd34933;
    data[ 192] =  'sd54120;
    data[ 193] =  'sd42272;
    data[ 194] =  'sd73754;
    data[ 195] =  'sd41599;
    data[ 196] =  'sd56929;
    data[ 197] = -'sd51344;
    data[ 198] =  'sd27128;
    data[ 199] =  'sd22836;
    data[ 200] =  'sd79377;
    data[ 201] =  'sd18333;
    data[ 202] = -'sd33198;
    data[ 203] = -'sd10745;
    data[ 204] =  'sd59057;
    data[ 205] =  'sd1856;
    data[ 206] =  'sd46400;
    data[ 207] =  'sd13113;
    data[ 208] =  'sd143;
    data[ 209] =  'sd3575;
    data[ 210] = -'sd74466;
    data[ 211] = -'sd59399;
    data[ 212] = -'sd10406;
    data[ 213] =  'sd67532;
    data[ 214] =  'sd49890;
    data[ 215] = -'sd63478;
    data[ 216] =  'sd51460;
    data[ 217] = -'sd24228;
    data[ 218] =  'sd49664;
    data[ 219] = -'sd69128;
    data[ 220] =  'sd74051;
    data[ 221] =  'sd49024;
    data[ 222] =  'sd78713;
    data[ 223] =  'sd1733;
    data[ 224] =  'sd43325;
    data[ 225] = -'sd63762;
    data[ 226] =  'sd44360;
    data[ 227] = -'sd37887;
    data[ 228] =  'sd35871;
    data[ 229] =  'sd77570;
    data[ 230] = -'sd26842;
    data[ 231] = -'sd15686;
    data[ 232] = -'sd64468;
    data[ 233] =  'sd26710;
    data[ 234] =  'sd12386;
    data[ 235] = -'sd18032;
    data[ 236] =  'sd40723;
    data[ 237] =  'sd35029;
    data[ 238] =  'sd56520;
    data[ 239] = -'sd61569;
    data[ 240] = -'sd64656;
    data[ 241] =  'sd22010;
    data[ 242] =  'sd58727;
    data[ 243] = -'sd6394;
    data[ 244] =  'sd3991;
    data[ 245] = -'sd64066;
    data[ 246] =  'sd36760;
    data[ 247] = -'sd64046;
    data[ 248] =  'sd37260;
    data[ 249] = -'sd51546;
    data[ 250] =  'sd22078;
    data[ 251] =  'sd60427;
    data[ 252] =  'sd36106;
    data[ 253] = -'sd80396;
    data[ 254] = -'sd43808;
    data[ 255] =  'sd51687;
    data[ 256] = -'sd18553;
    data[ 257] =  'sd27698;
    data[ 258] =  'sd37086;
    data[ 259] = -'sd55896;
    data[ 260] =  'sd77169;
    data[ 261] = -'sd36867;
    data[ 262] =  'sd61371;
    data[ 263] =  'sd59706;
    data[ 264] =  'sd18081;
    data[ 265] = -'sd39498;
    data[ 266] = -'sd4404;
    data[ 267] =  'sd53741;
    data[ 268] =  'sd32797;
    data[ 269] =  'sd720;
    data[ 270] =  'sd18000;
    data[ 271] = -'sd41523;
    data[ 272] = -'sd55029;
    data[ 273] = -'sd64997;
    data[ 274] =  'sd13485;
    data[ 275] =  'sd9443;
    data[ 276] =  'sd72234;
    data[ 277] =  'sd3599;
    data[ 278] = -'sd73866;
    data[ 279] = -'sd44399;
    data[ 280] =  'sd36912;
    data[ 281] = -'sd60246;
    data[ 282] = -'sd31581;
    data[ 283] =  'sd29680;
    data[ 284] = -'sd77205;
    data[ 285] =  'sd35967;
    data[ 286] =  'sd79970;
    data[ 287] =  'sd33158;
    data[ 288] =  'sd9745;
    data[ 289] =  'sd79784;
    data[ 290] =  'sd28508;
    data[ 291] =  'sd57336;
    data[ 292] = -'sd41169;
    data[ 293] = -'sd46179;
    data[ 294] = -'sd7588;
    data[ 295] = -'sd25859;
    data[ 296] =  'sd8889;
    data[ 297] =  'sd58384;
    data[ 298] = -'sd14969;
    data[ 299] = -'sd46543;
    data[ 300] = -'sd16688;
    data[ 301] =  'sd74323;
    data[ 302] =  'sd55824;
    data[ 303] = -'sd78969;
    data[ 304] = -'sd8133;
    data[ 305] = -'sd39484;
    data[ 306] = -'sd4054;
    data[ 307] =  'sd62491;
    data[ 308] = -'sd76135;
    data[ 309] =  'sd62717;
    data[ 310] = -'sd70485;
    data[ 311] =  'sd40126;
    data[ 312] =  'sd20104;
    data[ 313] =  'sd11077;
    data[ 314] = -'sd50757;
    data[ 315] =  'sd41803;
    data[ 316] =  'sd62029;
    data[ 317] =  'sd76156;
    data[ 318] = -'sd62192;
    data[ 319] = -'sd80231;
    data[ 320] = -'sd39683;
    data[ 321] = -'sd9029;
    data[ 322] = -'sd61884;
    data[ 323] = -'sd72531;
    data[ 324] = -'sd11024;
    data[ 325] =  'sd52082;
    data[ 326] = -'sd8678;
    data[ 327] = -'sd53109;
    data[ 328] = -'sd16997;
    data[ 329] =  'sd66598;
    data[ 330] =  'sd26540;
    data[ 331] =  'sd8136;
    data[ 332] =  'sd39559;
    data[ 333] =  'sd5929;
    data[ 334] = -'sd15616;
    data[ 335] = -'sd62718;
    data[ 336] =  'sd70460;
    data[ 337] = -'sd40751;
    data[ 338] = -'sd35729;
    data[ 339] = -'sd74020;
    data[ 340] = -'sd48249;
    data[ 341] = -'sd59338;
    data[ 342] = -'sd8881;
    data[ 343] = -'sd58184;
    data[ 344] =  'sd19969;
    data[ 345] =  'sd7702;
    data[ 346] =  'sd28709;
    data[ 347] =  'sd62361;
    data[ 348] = -'sd79385;
    data[ 349] = -'sd18533;
    data[ 350] =  'sd28198;
    data[ 351] =  'sd49586;
    data[ 352] = -'sd71078;
    data[ 353] =  'sd25301;
    data[ 354] = -'sd22839;
    data[ 355] = -'sd79452;
    data[ 356] = -'sd20208;
    data[ 357] = -'sd13677;
    data[ 358] = -'sd14243;
    data[ 359] = -'sd28393;
    data[ 360] = -'sd54461;
    data[ 361] = -'sd50797;
    data[ 362] =  'sd40803;
    data[ 363] =  'sd37029;
    data[ 364] = -'sd57321;
    data[ 365] =  'sd41544;
    data[ 366] =  'sd55554;
    data[ 367] =  'sd78122;
    data[ 368] = -'sd13042;
    data[ 369] =  'sd1632;
    data[ 370] =  'sd40800;
    data[ 371] =  'sd36954;
    data[ 372] = -'sd59196;
    data[ 373] = -'sd5331;
    data[ 374] =  'sd30566;
    data[ 375] = -'sd55055;
    data[ 376] = -'sd65647;
    data[ 377] = -'sd2765;
    data[ 378] = -'sd69125;
    data[ 379] =  'sd74126;
    data[ 380] =  'sd50899;
    data[ 381] = -'sd38253;
    data[ 382] =  'sd26721;
    data[ 383] =  'sd12661;
    data[ 384] = -'sd11157;
    data[ 385] =  'sd48757;
    data[ 386] =  'sd72038;
    data[ 387] = -'sd1301;
    data[ 388] = -'sd32525;
    data[ 389] =  'sd6080;
    data[ 390] = -'sd11841;
    data[ 391] =  'sd31657;
    data[ 392] = -'sd27780;
    data[ 393] = -'sd39136;
    data[ 394] =  'sd4646;
    data[ 395] = -'sd47691;
    data[ 396] = -'sd45388;
    data[ 397] =  'sd12187;
    data[ 398] = -'sd23007;
    data[ 399] =  'sd80189;
    data[ 400] =  'sd38633;
    data[ 401] = -'sd17221;
    data[ 402] =  'sd60998;
    data[ 403] =  'sd50381;
    data[ 404] = -'sd51203;
    data[ 405] =  'sd30653;
    data[ 406] = -'sd52880;
    data[ 407] = -'sd11272;
    data[ 408] =  'sd45882;
    data[ 409] =  'sd163;
    data[ 410] =  'sd4075;
    data[ 411] = -'sd61966;
    data[ 412] = -'sd74581;
    data[ 413] = -'sd62274;
    data[ 414] =  'sd81560;
    data[ 415] =  'sd72908;
    data[ 416] =  'sd20449;
    data[ 417] =  'sd19702;
    data[ 418] =  'sd1027;
    data[ 419] =  'sd25675;
    data[ 420] = -'sd13489;
    data[ 421] = -'sd9543;
    data[ 422] = -'sd74734;
    data[ 423] = -'sd66099;
    data[ 424] = -'sd14065;
    data[ 425] = -'sd23943;
    data[ 426] =  'sd56789;
    data[ 427] = -'sd54844;
    data[ 428] = -'sd60372;
    data[ 429] = -'sd34731;
    data[ 430] = -'sd49070;
    data[ 431] = -'sd79863;
    data[ 432] = -'sd30483;
    data[ 433] =  'sd57130;
    data[ 434] = -'sd46319;
    data[ 435] = -'sd11088;
    data[ 436] =  'sd50482;
    data[ 437] = -'sd48678;
    data[ 438] = -'sd70063;
    data[ 439] =  'sd50676;
    data[ 440] = -'sd43828;
    data[ 441] =  'sd51187;
    data[ 442] = -'sd31053;
    data[ 443] =  'sd42880;
    data[ 444] = -'sd74887;
    data[ 445] = -'sd69924;
    data[ 446] =  'sd54151;
    data[ 447] =  'sd43047;
    data[ 448] = -'sd70712;
    data[ 449] =  'sd34451;
    data[ 450] =  'sd42070;
    data[ 451] =  'sd68704;
    data[ 452] =  'sd79190;
    data[ 453] =  'sd13658;
    data[ 454] =  'sd13768;
    data[ 455] =  'sd16518;
    data[ 456] = -'sd78573;
    data[ 457] =  'sd1767;
    data[ 458] =  'sd44175;
    data[ 459] = -'sd42512;
    data[ 460] = -'sd79754;
    data[ 461] = -'sd27758;
    data[ 462] = -'sd38586;
    data[ 463] =  'sd18396;
    data[ 464] = -'sd31623;
    data[ 465] =  'sd28630;
    data[ 466] =  'sd60386;
    data[ 467] =  'sd35081;
    data[ 468] =  'sd57820;
    data[ 469] = -'sd29069;
    data[ 470] = -'sd71361;
    data[ 471] =  'sd18226;
    data[ 472] = -'sd35873;
    data[ 473] = -'sd77620;
    data[ 474] =  'sd25592;
    data[ 475] = -'sd15564;
    data[ 476] = -'sd61418;
    data[ 477] = -'sd60881;
    data[ 478] = -'sd47456;
    data[ 479] = -'sd39513;
    data[ 480] = -'sd4779;
    data[ 481] =  'sd44366;
    data[ 482] = -'sd37737;
    data[ 483] =  'sd39621;
    data[ 484] =  'sd7479;
    data[ 485] =  'sd23134;
    data[ 486] = -'sd77014;
    data[ 487] =  'sd40742;
    data[ 488] =  'sd35504;
    data[ 489] =  'sd68395;
    data[ 490] =  'sd71465;
    data[ 491] = -'sd15626;
    data[ 492] = -'sd62968;
    data[ 493] =  'sd64210;
    data[ 494] = -'sd33160;
    data[ 495] = -'sd9795;
    data[ 496] = -'sd81034;
    data[ 497] = -'sd59758;
    data[ 498] = -'sd19381;
    data[ 499] =  'sd6998;
    data[ 500] =  'sd11109;
    data[ 501] = -'sd49957;
    data[ 502] =  'sd61803;
    data[ 503] =  'sd70506;
    data[ 504] = -'sd39601;
    data[ 505] = -'sd6979;
    data[ 506] = -'sd10634;
    data[ 507] =  'sd61832;
    data[ 508] =  'sd71231;
    data[ 509] = -'sd21476;
    data[ 510] = -'sd45377;
    data[ 511] =  'sd12462;
    data[ 512] = -'sd16132;
    data[ 513] = -'sd75618;
    data[ 514] =  'sd75642;
    data[ 515] = -'sd75042;
    data[ 516] = -'sd73799;
    data[ 517] = -'sd42724;
    data[ 518] =  'sd78787;
    data[ 519] =  'sd3583;
    data[ 520] = -'sd74266;
    data[ 521] = -'sd54399;
    data[ 522] = -'sd49247;
    data[ 523] =  'sd79553;
    data[ 524] =  'sd22733;
    data[ 525] =  'sd76802;
    data[ 526] = -'sd46042;
    data[ 527] = -'sd4163;
    data[ 528] =  'sd59766;
    data[ 529] =  'sd19581;
    data[ 530] = -'sd1998;
    data[ 531] = -'sd49950;
    data[ 532] =  'sd61978;
    data[ 533] =  'sd74881;
    data[ 534] =  'sd69774;
    data[ 535] = -'sd57901;
    data[ 536] =  'sd27044;
    data[ 537] =  'sd20736;
    data[ 538] =  'sd26877;
    data[ 539] =  'sd16561;
    data[ 540] = -'sd77498;
    data[ 541] =  'sd28642;
    data[ 542] =  'sd60686;
    data[ 543] =  'sd42581;
    data[ 544] =  'sd81479;
    data[ 545] =  'sd70883;
    data[ 546] = -'sd30176;
    data[ 547] =  'sd64805;
    data[ 548] = -'sd18285;
    data[ 549] =  'sd34398;
    data[ 550] =  'sd40745;
    data[ 551] =  'sd35579;
    data[ 552] =  'sd70270;
    data[ 553] = -'sd45501;
    data[ 554] =  'sd9362;
    data[ 555] =  'sd70209;
    data[ 556] = -'sd47026;
    data[ 557] = -'sd28763;
    data[ 558] = -'sd63711;
    data[ 559] =  'sd45635;
    data[ 560] = -'sd6012;
    data[ 561] =  'sd13541;
    data[ 562] =  'sd10843;
    data[ 563] = -'sd56607;
    data[ 564] =  'sd59394;
    data[ 565] =  'sd10281;
    data[ 566] = -'sd70657;
    data[ 567] =  'sd35826;
    data[ 568] =  'sd76445;
    data[ 569] = -'sd54967;
    data[ 570] = -'sd63447;
    data[ 571] =  'sd52235;
    data[ 572] = -'sd4853;
    data[ 573] =  'sd42516;
    data[ 574] =  'sd79854;
    data[ 575] =  'sd30258;
    data[ 576] = -'sd62755;
    data[ 577] =  'sd69535;
    data[ 578] = -'sd63876;
    data[ 579] =  'sd41510;
    data[ 580] =  'sd54704;
    data[ 581] =  'sd56872;
    data[ 582] = -'sd52769;
    data[ 583] = -'sd8497;
    data[ 584] = -'sd48584;
    data[ 585] = -'sd67713;
    data[ 586] = -'sd54415;
    data[ 587] = -'sd49647;
    data[ 588] =  'sd69553;
    data[ 589] = -'sd63426;
    data[ 590] =  'sd52760;
    data[ 591] =  'sd8272;
    data[ 592] =  'sd42959;
    data[ 593] = -'sd72912;
    data[ 594] = -'sd20549;
    data[ 595] = -'sd22202;
    data[ 596] = -'sd63527;
    data[ 597] =  'sd50235;
    data[ 598] = -'sd54853;
    data[ 599] = -'sd60597;
    data[ 600] = -'sd40356;
    data[ 601] = -'sd25854;
    data[ 602] =  'sd9014;
    data[ 603] =  'sd61509;
    data[ 604] =  'sd63156;
    data[ 605] = -'sd59510;
    data[ 606] = -'sd13181;
    data[ 607] = -'sd1843;
    data[ 608] = -'sd46075;
    data[ 609] = -'sd4988;
    data[ 610] =  'sd39141;
    data[ 611] = -'sd4521;
    data[ 612] =  'sd50816;
    data[ 613] = -'sd40328;
    data[ 614] = -'sd25154;
    data[ 615] =  'sd26514;
    data[ 616] =  'sd7486;
    data[ 617] =  'sd23309;
    data[ 618] = -'sd72639;
    data[ 619] = -'sd13724;
    data[ 620] = -'sd15418;
    data[ 621] = -'sd57768;
    data[ 622] =  'sd30369;
    data[ 623] = -'sd59980;
    data[ 624] = -'sd24931;
    data[ 625] =  'sd32089;
    data[ 626] = -'sd16980;
    data[ 627] =  'sd67023;
    data[ 628] =  'sd37165;
    data[ 629] = -'sd53921;
    data[ 630] = -'sd37297;
    data[ 631] =  'sd50621;
    data[ 632] = -'sd45203;
    data[ 633] =  'sd16812;
    data[ 634] = -'sd71223;
    data[ 635] =  'sd21676;
    data[ 636] =  'sd50377;
    data[ 637] = -'sd51303;
    data[ 638] =  'sd28153;
    data[ 639] =  'sd48461;
    data[ 640] =  'sd64638;
    data[ 641] = -'sd22460;
    data[ 642] = -'sd69977;
    data[ 643] =  'sd52826;
    data[ 644] =  'sd9922;
    data[ 645] = -'sd79632;
    data[ 646] = -'sd24708;
    data[ 647] =  'sd37664;
    data[ 648] = -'sd41446;
    data[ 649] = -'sd53104;
    data[ 650] = -'sd16872;
    data[ 651] =  'sd69723;
    data[ 652] = -'sd59176;
    data[ 653] = -'sd4831;
    data[ 654] =  'sd43066;
    data[ 655] = -'sd70237;
    data[ 656] =  'sd46326;
    data[ 657] =  'sd11263;
    data[ 658] = -'sd46107;
    data[ 659] = -'sd5788;
    data[ 660] =  'sd19141;
    data[ 661] = -'sd12998;
    data[ 662] =  'sd2732;
    data[ 663] =  'sd68300;
    data[ 664] =  'sd69090;
    data[ 665] = -'sd75001;
    data[ 666] = -'sd72774;
    data[ 667] = -'sd17099;
    data[ 668] =  'sd64048;
    data[ 669] = -'sd37210;
    data[ 670] =  'sd52796;
    data[ 671] =  'sd9172;
    data[ 672] =  'sd65459;
    data[ 673] = -'sd1935;
    data[ 674] = -'sd48375;
    data[ 675] = -'sd62488;
    data[ 676] =  'sd76210;
    data[ 677] = -'sd60842;
    data[ 678] = -'sd46481;
    data[ 679] = -'sd15138;
    data[ 680] = -'sd50768;
    data[ 681] =  'sd41528;
    data[ 682] =  'sd55154;
    data[ 683] =  'sd68122;
    data[ 684] =  'sd64640;
    data[ 685] = -'sd22410;
    data[ 686] = -'sd68727;
    data[ 687] = -'sd79765;
    data[ 688] = -'sd28033;
    data[ 689] = -'sd45461;
    data[ 690] =  'sd10362;
    data[ 691] = -'sd68632;
    data[ 692] = -'sd77390;
    data[ 693] =  'sd31342;
    data[ 694] = -'sd35655;
    data[ 695] = -'sd72170;
    data[ 696] = -'sd1999;
    data[ 697] = -'sd49975;
    data[ 698] =  'sd61353;
    data[ 699] =  'sd59256;
    data[ 700] =  'sd6831;
    data[ 701] =  'sd6934;
    data[ 702] =  'sd9509;
    data[ 703] =  'sd73884;
    data[ 704] =  'sd44849;
    data[ 705] = -'sd25662;
    data[ 706] =  'sd13814;
    data[ 707] =  'sd17668;
    data[ 708] = -'sd49823;
    data[ 709] =  'sd65153;
    data[ 710] = -'sd9585;
    data[ 711] = -'sd75784;
    data[ 712] =  'sd71492;
    data[ 713] = -'sd14951;
    data[ 714] = -'sd46093;
    data[ 715] = -'sd5438;
    data[ 716] =  'sd27891;
    data[ 717] =  'sd41911;
    data[ 718] =  'sd64729;
    data[ 719] = -'sd20185;
    data[ 720] = -'sd13102;
    data[ 721] =  'sd132;
    data[ 722] =  'sd3300;
    data[ 723] = -'sd81341;
    data[ 724] = -'sd67433;
    data[ 725] = -'sd47415;
    data[ 726] = -'sd38488;
    data[ 727] =  'sd20846;
    data[ 728] =  'sd29627;
    data[ 729] = -'sd78530;
    data[ 730] =  'sd2842;
    data[ 731] =  'sd71050;
    data[ 732] = -'sd26001;
    data[ 733] =  'sd5339;
    data[ 734] = -'sd30366;
    data[ 735] =  'sd60055;
    data[ 736] =  'sd26806;
    data[ 737] =  'sd14786;
    data[ 738] =  'sd41968;
    data[ 739] =  'sd66154;
    data[ 740] =  'sd15440;
    data[ 741] =  'sd58318;
    data[ 742] = -'sd16619;
    data[ 743] =  'sd76048;
    data[ 744] = -'sd64892;
    data[ 745] =  'sd16110;
    data[ 746] =  'sd75068;
    data[ 747] =  'sd74449;
    data[ 748] =  'sd58974;
    data[ 749] = -'sd219;
    data[ 750] = -'sd5475;
    data[ 751] =  'sd26966;
    data[ 752] =  'sd18786;
    data[ 753] = -'sd21873;
    data[ 754] = -'sd55302;
    data[ 755] = -'sd71822;
    data[ 756] =  'sd6701;
    data[ 757] =  'sd3684;
    data[ 758] = -'sd71741;
    data[ 759] =  'sd8726;
    data[ 760] =  'sd54309;
    data[ 761] =  'sd46997;
    data[ 762] =  'sd28038;
    data[ 763] =  'sd45586;
    data[ 764] = -'sd7237;
    data[ 765] = -'sd17084;
    data[ 766] =  'sd64423;
    data[ 767] = -'sd27835;
    data[ 768] = -'sd40511;
    data[ 769] = -'sd29729;
    data[ 770] =  'sd75980;
    data[ 771] = -'sd66592;
    data[ 772] = -'sd26390;
    data[ 773] = -'sd4386;
    data[ 774] =  'sd54191;
    data[ 775] =  'sd44047;
    data[ 776] = -'sd45712;
    data[ 777] =  'sd4087;
    data[ 778] = -'sd61666;
    data[ 779] = -'sd67081;
    data[ 780] = -'sd38615;
    data[ 781] =  'sd17671;
    data[ 782] = -'sd49748;
    data[ 783] =  'sd67028;
    data[ 784] =  'sd37290;
    data[ 785] = -'sd50796;
    data[ 786] =  'sd40828;
    data[ 787] =  'sd37654;
    data[ 788] = -'sd41696;
    data[ 789] = -'sd59354;
    data[ 790] = -'sd9281;
    data[ 791] = -'sd68184;
    data[ 792] = -'sd66190;
    data[ 793] = -'sd16340;
    data[ 794] = -'sd80818;
    data[ 795] = -'sd54358;
    data[ 796] = -'sd48222;
    data[ 797] = -'sd58663;
    data[ 798] =  'sd7994;
    data[ 799] =  'sd36009;
    data[ 800] =  'sd81020;
    data[ 801] =  'sd59408;
    data[ 802] =  'sd10631;
    data[ 803] = -'sd61907;
    data[ 804] = -'sd73106;
    data[ 805] = -'sd25399;
    data[ 806] =  'sd20389;
    data[ 807] =  'sd18202;
    data[ 808] = -'sd36473;
    data[ 809] =  'sd71221;
    data[ 810] = -'sd21726;
    data[ 811] = -'sd51627;
    data[ 812] =  'sd20053;
    data[ 813] =  'sd9802;
    data[ 814] =  'sd81209;
    data[ 815] =  'sd64133;
    data[ 816] = -'sd35085;
    data[ 817] = -'sd57920;
    data[ 818] =  'sd26569;
    data[ 819] =  'sd8861;
    data[ 820] =  'sd57684;
    data[ 821] = -'sd32469;
    data[ 822] =  'sd7480;
    data[ 823] =  'sd23159;
    data[ 824] = -'sd76389;
    data[ 825] =  'sd56367;
    data[ 826] = -'sd65394;
    data[ 827] =  'sd3560;
    data[ 828] = -'sd74841;
    data[ 829] = -'sd68774;
    data[ 830] = -'sd80940;
    data[ 831] = -'sd57408;
    data[ 832] =  'sd39369;
    data[ 833] =  'sd1179;
    data[ 834] =  'sd29475;
    data[ 835] =  'sd81511;
    data[ 836] =  'sd71683;
    data[ 837] = -'sd10176;
    data[ 838] =  'sd73282;
    data[ 839] =  'sd29799;
    data[ 840] = -'sd74230;
    data[ 841] = -'sd53499;
    data[ 842] = -'sd26747;
    data[ 843] = -'sd13311;
    data[ 844] = -'sd5093;
    data[ 845] =  'sd36516;
    data[ 846] = -'sd70146;
    data[ 847] =  'sd48601;
    data[ 848] =  'sd68138;
    data[ 849] =  'sd65040;
    data[ 850] = -'sd12410;
    data[ 851] =  'sd17432;
    data[ 852] = -'sd55723;
    data[ 853] =  'sd81494;
    data[ 854] =  'sd71258;
    data[ 855] = -'sd20801;
    data[ 856] = -'sd28502;
    data[ 857] = -'sd57186;
    data[ 858] =  'sd44919;
    data[ 859] = -'sd23912;
    data[ 860] =  'sd57564;
    data[ 861] = -'sd35469;
    data[ 862] = -'sd67520;
    data[ 863] = -'sd49590;
    data[ 864] =  'sd70978;
    data[ 865] = -'sd27801;
    data[ 866] = -'sd39661;
    data[ 867] = -'sd8479;
    data[ 868] = -'sd48134;
    data[ 869] = -'sd56463;
    data[ 870] =  'sd62994;
    data[ 871] = -'sd63560;
    data[ 872] =  'sd49410;
    data[ 873] = -'sd75478;
    data[ 874] =  'sd79142;
    data[ 875] =  'sd12458;
    data[ 876] = -'sd16232;
    data[ 877] = -'sd78118;
    data[ 878] =  'sd13142;
    data[ 879] =  'sd868;
    data[ 880] =  'sd21700;
    data[ 881] =  'sd50977;
    data[ 882] = -'sd36303;
    data[ 883] =  'sd75471;
    data[ 884] = -'sd79317;
    data[ 885] = -'sd16833;
    data[ 886] =  'sd70698;
    data[ 887] = -'sd34801;
    data[ 888] = -'sd50820;
    data[ 889] =  'sd40228;
    data[ 890] =  'sd22654;
    data[ 891] =  'sd74827;
    data[ 892] =  'sd68424;
    data[ 893] =  'sd72190;
    data[ 894] =  'sd2499;
    data[ 895] =  'sd62475;
    data[ 896] = -'sd76535;
    data[ 897] =  'sd52717;
    data[ 898] =  'sd7197;
    data[ 899] =  'sd16084;
    data[ 900] =  'sd74418;
    data[ 901] =  'sd58199;
    data[ 902] = -'sd19594;
    data[ 903] =  'sd1673;
    data[ 904] =  'sd41825;
    data[ 905] =  'sd62579;
    data[ 906] = -'sd73935;
    data[ 907] = -'sd46124;
    data[ 908] = -'sd6213;
    data[ 909] =  'sd8516;
    data[ 910] =  'sd49059;
    data[ 911] =  'sd79588;
    data[ 912] =  'sd23608;
    data[ 913] = -'sd65164;
    data[ 914] =  'sd9310;
    data[ 915] =  'sd68909;
    data[ 916] = -'sd79526;
    data[ 917] = -'sd22058;
    data[ 918] = -'sd59927;
    data[ 919] = -'sd23606;
    data[ 920] =  'sd65214;
    data[ 921] = -'sd8060;
    data[ 922] = -'sd37659;
    data[ 923] =  'sd41571;
    data[ 924] =  'sd56229;
    data[ 925] = -'sd68844;
    data[ 926] =  'sd81151;
    data[ 927] =  'sd62683;
    data[ 928] = -'sd71335;
    data[ 929] =  'sd18876;
    data[ 930] = -'sd19623;
    data[ 931] =  'sd948;
    data[ 932] =  'sd23700;
    data[ 933] = -'sd62864;
    data[ 934] =  'sd66810;
    data[ 935] =  'sd31840;
    data[ 936] = -'sd23205;
    data[ 937] =  'sd75239;
    data[ 938] =  'sd78724;
    data[ 939] =  'sd2008;
    data[ 940] =  'sd50200;
    data[ 941] = -'sd55728;
    data[ 942] =  'sd81369;
    data[ 943] =  'sd68133;
    data[ 944] =  'sd64915;
    data[ 945] = -'sd15535;
    data[ 946] = -'sd60693;
    data[ 947] = -'sd42756;
    data[ 948] =  'sd77987;
    data[ 949] = -'sd16417;
    data[ 950] =  'sd81098;
    data[ 951] =  'sd61358;
    data[ 952] =  'sd59381;
    data[ 953] =  'sd9956;
    data[ 954] = -'sd78782;
    data[ 955] = -'sd3458;
    data[ 956] =  'sd77391;
    data[ 957] = -'sd31317;
    data[ 958] =  'sd36280;
    data[ 959] = -'sd76046;
    data[ 960] =  'sd64942;
    data[ 961] = -'sd14860;
    data[ 962] = -'sd43818;
    data[ 963] =  'sd51437;
    data[ 964] = -'sd24803;
    data[ 965] =  'sd35289;
    data[ 966] =  'sd63020;
    data[ 967] = -'sd62910;
    data[ 968] =  'sd65660;
    data[ 969] =  'sd3090;
    data[ 970] =  'sd77250;
    data[ 971] = -'sd34842;
    data[ 972] = -'sd51845;
    data[ 973] =  'sd14603;
    data[ 974] =  'sd37393;
    data[ 975] = -'sd48221;
    data[ 976] = -'sd58638;
    data[ 977] =  'sd8619;
    data[ 978] =  'sd51634;
    data[ 979] = -'sd19878;
    data[ 980] = -'sd5427;
    data[ 981] =  'sd28166;
    data[ 982] =  'sd48786;
    data[ 983] =  'sd72763;
    data[ 984] =  'sd16824;
    data[ 985] = -'sd70923;
    data[ 986] =  'sd29176;
    data[ 987] =  'sd74036;
    data[ 988] =  'sd48649;
    data[ 989] =  'sd69338;
    data[ 990] = -'sd68801;
    data[ 991] = -'sd81615;
    data[ 992] = -'sd74283;
    data[ 993] = -'sd54824;
    data[ 994] = -'sd59872;
    data[ 995] = -'sd22231;
    data[ 996] = -'sd64252;
    data[ 997] =  'sd32110;
    data[ 998] = -'sd16455;
    data[ 999] =  'sd80148;
    data[1000] =  'sd37608;
    data[1001] = -'sd42846;
    data[1002] =  'sd75737;
    data[1003] = -'sd72667;
    data[1004] = -'sd14424;
    data[1005] = -'sd32918;
    data[1006] = -'sd3745;
    data[1007] =  'sd70216;
    data[1008] = -'sd46851;
    data[1009] = -'sd24388;
    data[1010] =  'sd45664;
    data[1011] = -'sd5287;
    data[1012] =  'sd31666;
    data[1013] = -'sd27555;
    data[1014] = -'sd33511;
    data[1015] = -'sd18570;
    data[1016] =  'sd27273;
    data[1017] =  'sd26461;
    data[1018] =  'sd6161;
    data[1019] = -'sd9816;
    data[1020] = -'sd81559;
    data[1021] = -'sd72883;
    data[1022] = -'sd19824;
    data[1023] = -'sd4077;
    data[1024] =  'sd61916;
    data[1025] =  'sd73331;
    data[1026] =  'sd31024;
    data[1027] = -'sd43605;
    data[1028] =  'sd56762;
    data[1029] = -'sd55519;
    data[1030] = -'sd77247;
    data[1031] =  'sd34917;
    data[1032] =  'sd53720;
    data[1033] =  'sd32272;
    data[1034] = -'sd12405;
    data[1035] =  'sd17557;
    data[1036] = -'sd52598;
    data[1037] = -'sd4222;
    data[1038] =  'sd58291;
    data[1039] = -'sd17294;
    data[1040] =  'sd59173;
    data[1041] =  'sd4756;
    data[1042] = -'sd44941;
    data[1043] =  'sd23362;
    data[1044] = -'sd71314;
    data[1045] =  'sd19401;
    data[1046] = -'sd6498;
    data[1047] =  'sd1391;
    data[1048] =  'sd34775;
    data[1049] =  'sd50170;
    data[1050] = -'sd56478;
    data[1051] =  'sd62619;
    data[1052] = -'sd72935;
    data[1053] = -'sd21124;
    data[1054] = -'sd36577;
    data[1055] =  'sd68621;
    data[1056] =  'sd77115;
    data[1057] = -'sd38217;
    data[1058] =  'sd27621;
    data[1059] =  'sd35161;
    data[1060] =  'sd59820;
    data[1061] =  'sd20931;
    data[1062] =  'sd31752;
    data[1063] = -'sd25405;
    data[1064] =  'sd20239;
    data[1065] =  'sd14452;
    data[1066] =  'sd33618;
    data[1067] =  'sd21245;
    data[1068] =  'sd39602;
    data[1069] =  'sd7004;
    data[1070] =  'sd11259;
    data[1071] = -'sd46207;
    data[1072] = -'sd8288;
    data[1073] = -'sd43359;
    data[1074] =  'sd62912;
    data[1075] = -'sd65610;
    data[1076] = -'sd1840;
    data[1077] = -'sd46000;
    data[1078] = -'sd3113;
    data[1079] = -'sd77825;
    data[1080] =  'sd20467;
    data[1081] =  'sd20152;
    data[1082] =  'sd12277;
    data[1083] = -'sd20757;
    data[1084] = -'sd27402;
    data[1085] = -'sd29686;
    data[1086] =  'sd77055;
    data[1087] = -'sd39717;
    data[1088] = -'sd9879;
    data[1089] =  'sd80707;
    data[1090] =  'sd51583;
    data[1091] = -'sd21153;
    data[1092] = -'sd37302;
    data[1093] =  'sd50496;
    data[1094] = -'sd48328;
    data[1095] = -'sd61313;
    data[1096] = -'sd58256;
    data[1097] =  'sd18169;
    data[1098] = -'sd37298;
    data[1099] =  'sd50596;
    data[1100] = -'sd45828;
    data[1101] =  'sd1187;
    data[1102] =  'sd29675;
    data[1103] = -'sd77330;
    data[1104] =  'sd32842;
    data[1105] =  'sd1845;
    data[1106] =  'sd46125;
    data[1107] =  'sd6238;
    data[1108] = -'sd7891;
    data[1109] = -'sd33434;
    data[1110] = -'sd16645;
    data[1111] =  'sd75398;
    data[1112] = -'sd81142;
    data[1113] = -'sd62458;
    data[1114] =  'sd76960;
    data[1115] = -'sd42092;
    data[1116] = -'sd69254;
    data[1117] =  'sd70901;
    data[1118] = -'sd29726;
    data[1119] =  'sd76055;
    data[1120] = -'sd64717;
    data[1121] =  'sd20485;
    data[1122] =  'sd20602;
    data[1123] =  'sd23527;
    data[1124] = -'sd67189;
    data[1125] = -'sd41315;
    data[1126] = -'sd49829;
    data[1127] =  'sd65003;
    data[1128] = -'sd13335;
    data[1129] = -'sd5693;
    data[1130] =  'sd21516;
    data[1131] =  'sd46377;
    data[1132] =  'sd12538;
    data[1133] = -'sd14232;
    data[1134] = -'sd28118;
    data[1135] = -'sd47586;
    data[1136] = -'sd42763;
    data[1137] =  'sd77812;
    data[1138] = -'sd20792;
    data[1139] = -'sd28277;
    data[1140] = -'sd51561;
    data[1141] =  'sd21703;
    data[1142] =  'sd51052;
    data[1143] = -'sd34428;
    data[1144] = -'sd41495;
    data[1145] = -'sd54329;
    data[1146] = -'sd47497;
    data[1147] = -'sd40538;
    data[1148] = -'sd30404;
    data[1149] =  'sd59105;
    data[1150] =  'sd3056;
    data[1151] =  'sd76400;
    data[1152] = -'sd56092;
    data[1153] =  'sd72269;
    data[1154] =  'sd4474;
    data[1155] = -'sd51991;
    data[1156] =  'sd10953;
    data[1157] = -'sd53857;
    data[1158] = -'sd35697;
    data[1159] = -'sd73220;
    data[1160] = -'sd28249;
    data[1161] = -'sd50861;
    data[1162] =  'sd39203;
    data[1163] = -'sd2971;
    data[1164] = -'sd74275;
    data[1165] = -'sd54624;
    data[1166] = -'sd54872;
    data[1167] = -'sd61072;
    data[1168] = -'sd52231;
    data[1169] =  'sd4953;
    data[1170] = -'sd40016;
    data[1171] = -'sd17354;
    data[1172] =  'sd57673;
    data[1173] = -'sd32744;
    data[1174] =  'sd605;
    data[1175] =  'sd15125;
    data[1176] =  'sd50443;
    data[1177] = -'sd49653;
    data[1178] =  'sd69403;
    data[1179] = -'sd67176;
    data[1180] = -'sd40990;
    data[1181] = -'sd41704;
    data[1182] = -'sd59554;
    data[1183] = -'sd14281;
    data[1184] = -'sd29343;
    data[1185] = -'sd78211;
    data[1186] =  'sd10817;
    data[1187] = -'sd57257;
    data[1188] =  'sd43144;
    data[1189] = -'sd68287;
    data[1190] = -'sd68765;
    data[1191] = -'sd80715;
    data[1192] = -'sd51783;
    data[1193] =  'sd16153;
    data[1194] =  'sd76143;
    data[1195] = -'sd62517;
    data[1196] =  'sd75485;
    data[1197] = -'sd78967;
    data[1198] = -'sd8083;
    data[1199] = -'sd38234;
    data[1200] =  'sd27196;
    data[1201] =  'sd24536;
    data[1202] = -'sd41964;
    data[1203] = -'sd66054;
    data[1204] = -'sd12940;
    data[1205] =  'sd4182;
    data[1206] = -'sd59291;
    data[1207] = -'sd7706;
    data[1208] = -'sd28809;
    data[1209] = -'sd64861;
    data[1210] =  'sd16885;
    data[1211] = -'sd69398;
    data[1212] =  'sd67301;
    data[1213] =  'sd44115;
    data[1214] = -'sd44012;
    data[1215] =  'sd46587;
    data[1216] =  'sd17788;
    data[1217] = -'sd46823;
    data[1218] = -'sd23688;
    data[1219] =  'sd63164;
    data[1220] = -'sd59310;
    data[1221] = -'sd8181;
    data[1222] = -'sd40684;
    data[1223] = -'sd34054;
    data[1224] = -'sd32145;
    data[1225] =  'sd15580;
    data[1226] =  'sd61818;
    data[1227] =  'sd70881;
    data[1228] = -'sd30226;
    data[1229] =  'sd63555;
    data[1230] = -'sd49535;
    data[1231] =  'sd72353;
    data[1232] =  'sd6574;
    data[1233] =  'sd509;
    data[1234] =  'sd12725;
    data[1235] = -'sd9557;
    data[1236] = -'sd75084;
    data[1237] = -'sd74849;
    data[1238] = -'sd68974;
    data[1239] =  'sd77901;
    data[1240] = -'sd18567;
    data[1241] =  'sd27348;
    data[1242] =  'sd28336;
    data[1243] =  'sd53036;
    data[1244] =  'sd15172;
    data[1245] =  'sd51618;
    data[1246] = -'sd20278;
    data[1247] = -'sd15427;
    data[1248] = -'sd57993;
    data[1249] =  'sd24744;
    data[1250] = -'sd36764;
    data[1251] =  'sd63946;
    data[1252] = -'sd39760;
    data[1253] = -'sd10954;
    data[1254] =  'sd53832;
    data[1255] =  'sd35072;
    data[1256] =  'sd57595;
    data[1257] = -'sd34694;
    data[1258] = -'sd48145;
    data[1259] = -'sd56738;
    data[1260] =  'sd56119;
    data[1261] = -'sd71594;
    data[1262] =  'sd12401;
    data[1263] = -'sd17657;
    data[1264] =  'sd50098;
    data[1265] = -'sd58278;
    data[1266] =  'sd17619;
    data[1267] = -'sd51048;
    data[1268] =  'sd34528;
    data[1269] =  'sd43995;
    data[1270] = -'sd47012;
    data[1271] = -'sd28413;
    data[1272] = -'sd54961;
    data[1273] = -'sd63297;
    data[1274] =  'sd55985;
    data[1275] = -'sd74944;
    data[1276] = -'sd71349;
    data[1277] =  'sd18526;
    data[1278] = -'sd28373;
    data[1279] = -'sd53961;
    data[1280] = -'sd38297;
    data[1281] =  'sd25621;
    data[1282] = -'sd14839;
    data[1283] = -'sd43293;
    data[1284] =  'sd64562;
    data[1285] = -'sd24360;
    data[1286] =  'sd46364;
    data[1287] =  'sd12213;
    data[1288] = -'sd22357;
    data[1289] = -'sd67402;
    data[1290] = -'sd46640;
    data[1291] = -'sd19113;
    data[1292] =  'sd13698;
    data[1293] =  'sd14768;
    data[1294] =  'sd41518;
    data[1295] =  'sd54904;
    data[1296] =  'sd61872;
    data[1297] =  'sd72231;
    data[1298] =  'sd3524;
    data[1299] = -'sd75741;
    data[1300] =  'sd72567;
    data[1301] =  'sd11924;
    data[1302] = -'sd29582;
    data[1303] =  'sd79655;
    data[1304] =  'sd25283;
    data[1305] = -'sd23289;
    data[1306] =  'sd73139;
    data[1307] =  'sd26224;
    data[1308] =  'sd236;
    data[1309] =  'sd5900;
    data[1310] = -'sd16341;
    data[1311] = -'sd80843;
    data[1312] = -'sd54983;
    data[1313] = -'sd63847;
    data[1314] =  'sd42235;
    data[1315] =  'sd72829;
    data[1316] =  'sd18474;
    data[1317] = -'sd29673;
    data[1318] =  'sd77380;
    data[1319] = -'sd31592;
    data[1320] =  'sd29405;
    data[1321] =  'sd79761;
    data[1322] =  'sd27933;
    data[1323] =  'sd42961;
    data[1324] = -'sd72862;
    data[1325] = -'sd19299;
    data[1326] =  'sd9048;
    data[1327] =  'sd62359;
    data[1328] = -'sd79435;
    data[1329] = -'sd19783;
    data[1330] = -'sd3052;
    data[1331] = -'sd76300;
    data[1332] =  'sd58592;
    data[1333] = -'sd9769;
    data[1334] = -'sd80384;
    data[1335] = -'sd43508;
    data[1336] =  'sd59187;
    data[1337] =  'sd5106;
    data[1338] = -'sd36191;
    data[1339] =  'sd78271;
    data[1340] = -'sd9317;
    data[1341] = -'sd69084;
    data[1342] =  'sd75151;
    data[1343] =  'sd76524;
    data[1344] = -'sd52992;
    data[1345] = -'sd14072;
    data[1346] = -'sd24118;
    data[1347] =  'sd52414;
    data[1348] = -'sd378;
    data[1349] = -'sd9450;
    data[1350] = -'sd72409;
    data[1351] = -'sd7974;
    data[1352] = -'sd35509;
    data[1353] = -'sd68520;
    data[1354] = -'sd74590;
    data[1355] = -'sd62499;
    data[1356] =  'sd75935;
    data[1357] = -'sd67717;
    data[1358] = -'sd54515;
    data[1359] = -'sd52147;
    data[1360] =  'sd7053;
    data[1361] =  'sd12484;
    data[1362] = -'sd15582;
    data[1363] = -'sd61868;
    data[1364] = -'sd72131;
    data[1365] = -'sd1024;
    data[1366] = -'sd25600;
    data[1367] =  'sd15364;
    data[1368] =  'sd56418;
    data[1369] = -'sd64119;
    data[1370] =  'sd35435;
    data[1371] =  'sd66670;
    data[1372] =  'sd28340;
    data[1373] =  'sd53136;
    data[1374] =  'sd17672;
    data[1375] = -'sd49723;
    data[1376] =  'sd67653;
    data[1377] =  'sd52915;
    data[1378] =  'sd12147;
    data[1379] = -'sd24007;
    data[1380] =  'sd55189;
    data[1381] =  'sd68997;
    data[1382] = -'sd77326;
    data[1383] =  'sd32942;
    data[1384] =  'sd4345;
    data[1385] = -'sd55216;
    data[1386] = -'sd69672;
    data[1387] =  'sd60451;
    data[1388] =  'sd36706;
    data[1389] = -'sd65396;
    data[1390] =  'sd3510;
    data[1391] = -'sd76091;
    data[1392] =  'sd63817;
    data[1393] = -'sd42985;
    data[1394] =  'sd72262;
    data[1395] =  'sd4299;
    data[1396] = -'sd56366;
    data[1397] =  'sd65419;
    data[1398] = -'sd2935;
    data[1399] = -'sd73375;
    data[1400] = -'sd32124;
    data[1401] =  'sd16105;
    data[1402] =  'sd74943;
    data[1403] =  'sd71324;
    data[1404] = -'sd19151;
    data[1405] =  'sd12748;
    data[1406] = -'sd8982;
    data[1407] = -'sd60709;
    data[1408] = -'sd43156;
    data[1409] =  'sd67987;
    data[1410] =  'sd61265;
    data[1411] =  'sd57056;
    data[1412] = -'sd48169;
    data[1413] = -'sd57338;
    data[1414] =  'sd41119;
    data[1415] =  'sd44929;
    data[1416] = -'sd23662;
    data[1417] =  'sd63814;
    data[1418] = -'sd43060;
    data[1419] =  'sd70387;
    data[1420] = -'sd42576;
    data[1421] = -'sd81354;
    data[1422] = -'sd67758;
    data[1423] = -'sd55540;
    data[1424] = -'sd77772;
    data[1425] =  'sd21792;
    data[1426] =  'sd53277;
    data[1427] =  'sd21197;
    data[1428] =  'sd38402;
    data[1429] = -'sd22996;
    data[1430] =  'sd80464;
    data[1431] =  'sd45508;
    data[1432] = -'sd9187;
    data[1433] = -'sd65834;
    data[1434] = -'sd7440;
    data[1435] = -'sd22159;
    data[1436] = -'sd62452;
    data[1437] =  'sd77110;
    data[1438] = -'sd38342;
    data[1439] =  'sd24496;
    data[1440] = -'sd42964;
    data[1441] =  'sd72787;
    data[1442] =  'sd17424;
    data[1443] = -'sd55923;
    data[1444] =  'sd76494;
    data[1445] = -'sd53742;
    data[1446] = -'sd32822;
    data[1447] = -'sd1345;
    data[1448] = -'sd33625;
    data[1449] = -'sd21420;
    data[1450] = -'sd43977;
    data[1451] =  'sd47462;
    data[1452] =  'sd39663;
    data[1453] =  'sd8529;
    data[1454] =  'sd49384;
    data[1455] = -'sd76128;
    data[1456] =  'sd62892;
    data[1457] = -'sd66110;
    data[1458] = -'sd14340;
    data[1459] = -'sd30818;
    data[1460] =  'sd48755;
    data[1461] =  'sd71988;
    data[1462] = -'sd2551;
    data[1463] = -'sd63775;
    data[1464] =  'sd44035;
    data[1465] = -'sd46012;
    data[1466] = -'sd3413;
    data[1467] =  'sd78516;
    data[1468] = -'sd3192;
    data[1469] = -'sd79800;
    data[1470] = -'sd28908;
    data[1471] = -'sd67336;
    data[1472] = -'sd44990;
    data[1473] =  'sd22137;
    data[1474] =  'sd61902;
    data[1475] =  'sd72981;
    data[1476] =  'sd22274;
    data[1477] =  'sd65327;
    data[1478] = -'sd5235;
    data[1479] =  'sd32966;
    data[1480] =  'sd4945;
    data[1481] = -'sd40216;
    data[1482] = -'sd22354;
    data[1483] = -'sd67327;
    data[1484] = -'sd44765;
    data[1485] =  'sd27762;
    data[1486] =  'sd38686;
    data[1487] = -'sd15896;
    data[1488] = -'sd69718;
    data[1489] =  'sd59301;
    data[1490] =  'sd7956;
    data[1491] =  'sd35059;
    data[1492] =  'sd57270;
    data[1493] = -'sd42819;
    data[1494] =  'sd76412;
    data[1495] = -'sd55792;
    data[1496] =  'sd79769;
    data[1497] =  'sd28133;
    data[1498] =  'sd47961;
    data[1499] =  'sd52138;
    data[1500] = -'sd7278;
    data[1501] = -'sd18109;
    data[1502] =  'sd38798;
    data[1503] = -'sd13096;
    data[1504] =  'sd282;
    data[1505] =  'sd7050;
    data[1506] =  'sd12409;
    data[1507] = -'sd17457;
    data[1508] =  'sd55098;
    data[1509] =  'sd66722;
    data[1510] =  'sd29640;
    data[1511] = -'sd78205;
    data[1512] =  'sd10967;
    data[1513] = -'sd53507;
    data[1514] = -'sd26947;
    data[1515] = -'sd18311;
    data[1516] =  'sd33748;
    data[1517] =  'sd24495;
    data[1518] = -'sd42989;
    data[1519] =  'sd72162;
    data[1520] =  'sd1799;
    data[1521] =  'sd44975;
    data[1522] = -'sd22512;
    data[1523] = -'sd71277;
    data[1524] =  'sd20326;
    data[1525] =  'sd16627;
    data[1526] = -'sd75848;
    data[1527] =  'sd69892;
    data[1528] = -'sd54951;
    data[1529] = -'sd63047;
    data[1530] =  'sd62235;
    data[1531] =  'sd81306;
    data[1532] =  'sd66558;
    data[1533] =  'sd25540;
    data[1534] = -'sd16864;
    data[1535] =  'sd69923;
    data[1536] = -'sd54176;
    data[1537] = -'sd43672;
    data[1538] =  'sd55087;
    data[1539] =  'sd66447;
    data[1540] =  'sd22765;
    data[1541] =  'sd77602;
    data[1542] = -'sd26042;
    data[1543] =  'sd4314;
    data[1544] = -'sd55991;
    data[1545] =  'sd74794;
    data[1546] =  'sd67599;
    data[1547] =  'sd51565;
    data[1548] = -'sd21603;
    data[1549] = -'sd48552;
    data[1550] = -'sd66913;
    data[1551] = -'sd34415;
    data[1552] = -'sd41170;
    data[1553] = -'sd46204;
    data[1554] = -'sd8213;
    data[1555] = -'sd41484;
    data[1556] = -'sd54054;
    data[1557] = -'sd40622;
    data[1558] = -'sd32504;
    data[1559] =  'sd6605;
    data[1560] =  'sd1284;
    data[1561] =  'sd32100;
    data[1562] = -'sd16705;
    data[1563] =  'sd73898;
    data[1564] =  'sd45199;
    data[1565] = -'sd16912;
    data[1566] =  'sd68723;
    data[1567] =  'sd79665;
    data[1568] =  'sd25533;
    data[1569] = -'sd17039;
    data[1570] =  'sd65548;
    data[1571] =  'sd290;
    data[1572] =  'sd7250;
    data[1573] =  'sd17409;
    data[1574] = -'sd56298;
    data[1575] =  'sd67119;
    data[1576] =  'sd39565;
    data[1577] =  'sd6079;
    data[1578] = -'sd11866;
    data[1579] =  'sd31032;
    data[1580] = -'sd43405;
    data[1581] =  'sd61762;
    data[1582] =  'sd69481;
    data[1583] = -'sd65226;
    data[1584] =  'sd7760;
    data[1585] =  'sd30159;
    data[1586] = -'sd65230;
    data[1587] =  'sd7660;
    data[1588] =  'sd27659;
    data[1589] =  'sd36111;
    data[1590] = -'sd80271;
    data[1591] = -'sd40683;
    data[1592] = -'sd34029;
    data[1593] = -'sd31520;
    data[1594] =  'sd31205;
    data[1595] = -'sd39080;
    data[1596] =  'sd6046;
    data[1597] = -'sd12691;
    data[1598] =  'sd10407;
    data[1599] = -'sd67507;
    data[1600] = -'sd49265;
    data[1601] =  'sd79103;
    data[1602] =  'sd11483;
    data[1603] = -'sd40607;
    data[1604] = -'sd32129;
    data[1605] =  'sd15980;
    data[1606] =  'sd71818;
    data[1607] = -'sd6801;
    data[1608] = -'sd6184;
    data[1609] =  'sd9241;
    data[1610] =  'sd67184;
    data[1611] =  'sd41190;
    data[1612] =  'sd46704;
    data[1613] =  'sd20713;
    data[1614] =  'sd26302;
    data[1615] =  'sd2186;
    data[1616] =  'sd54650;
    data[1617] =  'sd55522;
    data[1618] =  'sd77322;
    data[1619] = -'sd33042;
    data[1620] = -'sd6845;
    data[1621] = -'sd7284;
    data[1622] = -'sd18259;
    data[1623] =  'sd35048;
    data[1624] =  'sd56995;
    data[1625] = -'sd49694;
    data[1626] =  'sd68378;
    data[1627] =  'sd71040;
    data[1628] = -'sd26251;
    data[1629] = -'sd911;
    data[1630] = -'sd22775;
    data[1631] = -'sd77852;
    data[1632] =  'sd19792;
    data[1633] =  'sd3277;
    data[1634] = -'sd81916;
    data[1635] = -'sd81808;
    data[1636] = -'sd79108;
    data[1637] = -'sd11608;
    data[1638] =  'sd37482;
    data[1639] = -'sd45996;
    data[1640] = -'sd3013;
    data[1641] = -'sd75325;
    data[1642] = -'sd80874;
    data[1643] = -'sd55758;
    data[1644] =  'sd80619;
    data[1645] =  'sd49383;
    data[1646] = -'sd76153;
    data[1647] =  'sd62267;
    data[1648] = -'sd81735;
    data[1649] = -'sd77283;
    data[1650] =  'sd34017;
    data[1651] =  'sd31220;
    data[1652] = -'sd38705;
    data[1653] =  'sd15421;
    data[1654] =  'sd57843;
    data[1655] = -'sd28494;
    data[1656] = -'sd56986;
    data[1657] =  'sd49919;
    data[1658] = -'sd62753;
    data[1659] =  'sd69585;
    data[1660] = -'sd62626;
    data[1661] =  'sd72760;
    data[1662] =  'sd16749;
    data[1663] = -'sd72798;
    data[1664] = -'sd17699;
    data[1665] =  'sd49048;
    data[1666] =  'sd79313;
    data[1667] =  'sd16733;
    data[1668] = -'sd73198;
    data[1669] = -'sd27699;
    data[1670] = -'sd37111;
    data[1671] =  'sd55271;
    data[1672] =  'sd71047;
    data[1673] = -'sd26076;
    data[1674] =  'sd3464;
    data[1675] = -'sd77241;
    data[1676] =  'sd35067;
    data[1677] =  'sd57470;
    data[1678] = -'sd37819;
    data[1679] =  'sd37571;
    data[1680] = -'sd43771;
    data[1681] =  'sd52612;
    data[1682] =  'sd4572;
    data[1683] = -'sd49541;
    data[1684] =  'sd72203;
    data[1685] =  'sd2824;
    data[1686] =  'sd70600;
    data[1687] = -'sd37251;
    data[1688] =  'sd51771;
    data[1689] = -'sd16453;
    data[1690] =  'sd80198;
    data[1691] =  'sd38858;
    data[1692] = -'sd11596;
    data[1693] =  'sd37782;
    data[1694] = -'sd38496;
    data[1695] =  'sd20646;
    data[1696] =  'sd24627;
    data[1697] = -'sd39689;
    data[1698] = -'sd9179;
    data[1699] = -'sd65634;
    data[1700] = -'sd2440;
    data[1701] = -'sd61000;
    data[1702] = -'sd50431;
    data[1703] =  'sd49953;
    data[1704] = -'sd61903;
    data[1705] = -'sd73006;
    data[1706] = -'sd22899;
    data[1707] = -'sd80952;
    data[1708] = -'sd57708;
    data[1709] =  'sd31869;
    data[1710] = -'sd22480;
    data[1711] = -'sd70477;
    data[1712] =  'sd40326;
    data[1713] =  'sd25104;
    data[1714] = -'sd27764;
    data[1715] = -'sd38736;
    data[1716] =  'sd14646;
    data[1717] =  'sd38468;
    data[1718] = -'sd21346;
    data[1719] = -'sd42127;
    data[1720] = -'sd70129;
    data[1721] =  'sd49026;
    data[1722] =  'sd78763;
    data[1723] =  'sd2983;
    data[1724] =  'sd74575;
    data[1725] =  'sd62124;
    data[1726] =  'sd78531;
    data[1727] = -'sd2817;
    data[1728] = -'sd70425;
    data[1729] =  'sd41626;
    data[1730] =  'sd57604;
    data[1731] = -'sd34469;
    data[1732] = -'sd42520;
    data[1733] = -'sd79954;
    data[1734] = -'sd32758;
    data[1735] =  'sd255;
    data[1736] =  'sd6375;
    data[1737] = -'sd4466;
    data[1738] =  'sd52191;
    data[1739] = -'sd5953;
    data[1740] =  'sd15016;
    data[1741] =  'sd47718;
    data[1742] =  'sd46063;
    data[1743] =  'sd4688;
    data[1744] = -'sd46641;
    data[1745] = -'sd19138;
    data[1746] =  'sd13073;
    data[1747] = -'sd857;
    data[1748] = -'sd21425;
    data[1749] = -'sd44102;
    data[1750] =  'sd44337;
    data[1751] = -'sd38462;
    data[1752] =  'sd21496;
    data[1753] =  'sd45877;
    data[1754] =  'sd38;
    data[1755] =  'sd950;
    data[1756] =  'sd23750;
    data[1757] = -'sd61614;
    data[1758] = -'sd65781;
    data[1759] = -'sd6115;
    data[1760] =  'sd10966;
    data[1761] = -'sd53532;
    data[1762] = -'sd27572;
    data[1763] = -'sd33936;
    data[1764] = -'sd29195;
    data[1765] = -'sd74511;
    data[1766] = -'sd60524;
    data[1767] = -'sd38531;
    data[1768] =  'sd19771;
    data[1769] =  'sd2752;
    data[1770] =  'sd68800;
    data[1771] =  'sd81590;
    data[1772] =  'sd73658;
    data[1773] =  'sd39199;
    data[1774] = -'sd3071;
    data[1775] = -'sd76775;
    data[1776] =  'sd46717;
    data[1777] =  'sd21038;
    data[1778] =  'sd34427;
    data[1779] =  'sd41470;
    data[1780] =  'sd53704;
    data[1781] =  'sd31872;
    data[1782] = -'sd22405;
    data[1783] = -'sd68602;
    data[1784] = -'sd76640;
    data[1785] =  'sd50092;
    data[1786] = -'sd58428;
    data[1787] =  'sd13869;
    data[1788] =  'sd19043;
    data[1789] = -'sd15448;
    data[1790] = -'sd58518;
    data[1791] =  'sd11619;
    data[1792] = -'sd37207;
    data[1793] =  'sd52871;
    data[1794] =  'sd11047;
    data[1795] = -'sd51507;
    data[1796] =  'sd23053;
    data[1797] = -'sd79039;
    data[1798] = -'sd9883;
    data[1799] =  'sd80607;
    data[1800] =  'sd49083;
    data[1801] =  'sd80188;
    data[1802] =  'sd38608;
    data[1803] = -'sd17846;
    data[1804] =  'sd45373;
    data[1805] = -'sd12562;
    data[1806] =  'sd13632;
    data[1807] =  'sd13118;
    data[1808] =  'sd268;
    data[1809] =  'sd6700;
    data[1810] =  'sd3659;
    data[1811] = -'sd72366;
    data[1812] = -'sd6899;
    data[1813] = -'sd8634;
    data[1814] = -'sd52009;
    data[1815] =  'sd10503;
    data[1816] = -'sd65107;
    data[1817] =  'sd10735;
    data[1818] = -'sd59307;
    data[1819] = -'sd8106;
    data[1820] = -'sd38809;
    data[1821] =  'sd12821;
    data[1822] = -'sd7157;
    data[1823] = -'sd15084;
    data[1824] = -'sd49418;
    data[1825] =  'sd75278;
    data[1826] =  'sd79699;
    data[1827] =  'sd26383;
    data[1828] =  'sd4211;
    data[1829] = -'sd58566;
    data[1830] =  'sd10419;
    data[1831] = -'sd67207;
    data[1832] = -'sd41765;
    data[1833] = -'sd61079;
    data[1834] = -'sd52406;
    data[1835] =  'sd578;
    data[1836] =  'sd14450;
    data[1837] =  'sd33568;
    data[1838] =  'sd19995;
    data[1839] =  'sd8352;
    data[1840] =  'sd44959;
    data[1841] = -'sd22912;
    data[1842] = -'sd81277;
    data[1843] = -'sd65833;
    data[1844] = -'sd7415;
    data[1845] = -'sd21534;
    data[1846] = -'sd46827;
    data[1847] = -'sd23788;
    data[1848] =  'sd60664;
    data[1849] =  'sd42031;
    data[1850] =  'sd67729;
    data[1851] =  'sd54815;
    data[1852] =  'sd59647;
    data[1853] =  'sd16606;
    data[1854] = -'sd76373;
    data[1855] =  'sd56767;
    data[1856] = -'sd55394;
    data[1857] = -'sd74122;
    data[1858] = -'sd50799;
    data[1859] =  'sd40753;
    data[1860] =  'sd35779;
    data[1861] =  'sd75270;
    data[1862] =  'sd79499;
    data[1863] =  'sd21383;
    data[1864] =  'sd43052;
    data[1865] = -'sd70587;
    data[1866] =  'sd37576;
    data[1867] = -'sd43646;
    data[1868] =  'sd55737;
    data[1869] = -'sd81144;
    data[1870] = -'sd62508;
    data[1871] =  'sd75710;
    data[1872] = -'sd73342;
    data[1873] = -'sd31299;
    data[1874] =  'sd36730;
    data[1875] = -'sd64796;
    data[1876] =  'sd18510;
    data[1877] = -'sd28773;
    data[1878] = -'sd63961;
    data[1879] =  'sd39385;
    data[1880] =  'sd1579;
    data[1881] =  'sd39475;
    data[1882] =  'sd3829;
    data[1883] = -'sd68116;
    data[1884] = -'sd64490;
    data[1885] =  'sd26160;
    data[1886] = -'sd1364;
    data[1887] = -'sd34100;
    data[1888] = -'sd33295;
    data[1889] = -'sd13170;
    data[1890] = -'sd1568;
    data[1891] = -'sd39200;
    data[1892] =  'sd3046;
    data[1893] =  'sd76150;
    data[1894] = -'sd62342;
    data[1895] =  'sd79860;
    data[1896] =  'sd30408;
    data[1897] = -'sd59005;
    data[1898] = -'sd556;
    data[1899] = -'sd13900;
    data[1900] = -'sd19818;
    data[1901] = -'sd3927;
    data[1902] =  'sd65666;
    data[1903] =  'sd3240;
    data[1904] =  'sd81000;
    data[1905] =  'sd58908;
    data[1906] = -'sd1869;
    data[1907] = -'sd46725;
    data[1908] = -'sd21238;
    data[1909] = -'sd39427;
    data[1910] = -'sd2629;
    data[1911] = -'sd65725;
    data[1912] = -'sd4715;
    data[1913] =  'sd45966;
    data[1914] =  'sd2263;
    data[1915] =  'sd56575;
    data[1916] = -'sd60194;
    data[1917] = -'sd30281;
    data[1918] =  'sd62180;
    data[1919] =  'sd79931;
    data[1920] =  'sd32183;
    data[1921] = -'sd14630;
    data[1922] = -'sd38068;
    data[1923] =  'sd31346;
    data[1924] = -'sd35555;
    data[1925] = -'sd69670;
    data[1926] =  'sd60501;
    data[1927] =  'sd37956;
    data[1928] = -'sd34146;
    data[1929] = -'sd34445;
    data[1930] = -'sd41920;
    data[1931] = -'sd64954;
    data[1932] =  'sd14560;
    data[1933] =  'sd36318;
    data[1934] = -'sd75096;
    data[1935] = -'sd75149;
    data[1936] = -'sd76474;
    data[1937] =  'sd54242;
    data[1938] =  'sd45322;
    data[1939] = -'sd13837;
    data[1940] = -'sd18243;
    data[1941] =  'sd35448;
    data[1942] =  'sd66995;
    data[1943] =  'sd36465;
    data[1944] = -'sd71421;
    data[1945] =  'sd16726;
    data[1946] = -'sd73373;
    data[1947] = -'sd32074;
    data[1948] =  'sd17355;
    data[1949] = -'sd57648;
    data[1950] =  'sd33369;
    data[1951] =  'sd15020;
    data[1952] =  'sd47818;
    data[1953] =  'sd48563;
    data[1954] =  'sd67188;
    data[1955] =  'sd41290;
    data[1956] =  'sd49204;
    data[1957] = -'sd80628;
    data[1958] = -'sd49608;
    data[1959] =  'sd70528;
    data[1960] = -'sd39051;
    data[1961] =  'sd6771;
    data[1962] =  'sd5434;
    data[1963] = -'sd27991;
    data[1964] = -'sd44411;
    data[1965] =  'sd36612;
    data[1966] = -'sd67746;
    data[1967] = -'sd55240;
    data[1968] = -'sd70272;
    data[1969] =  'sd45451;
    data[1970] = -'sd10612;
    data[1971] =  'sd62382;
    data[1972] = -'sd78860;
    data[1973] = -'sd5408;
    data[1974] =  'sd28641;
    data[1975] =  'sd60661;
    data[1976] =  'sd41956;
    data[1977] =  'sd65854;
    data[1978] =  'sd7940;
    data[1979] =  'sd34659;
    data[1980] =  'sd47270;
    data[1981] =  'sd34863;
    data[1982] =  'sd52370;
    data[1983] = -'sd1478;
    data[1984] = -'sd36950;
    data[1985] =  'sd59296;
    data[1986] =  'sd7831;
    data[1987] =  'sd31934;
    data[1988] = -'sd20855;
    data[1989] = -'sd29852;
    data[1990] =  'sd72905;
    data[1991] =  'sd20374;
    data[1992] =  'sd17827;
    data[1993] = -'sd45848;
    data[1994] =  'sd687;
    data[1995] =  'sd17175;
    data[1996] = -'sd62148;
    data[1997] = -'sd79131;
    data[1998] = -'sd12183;
    data[1999] =  'sd23107;
    data[2000] = -'sd77689;
    data[2001] =  'sd23867;
    data[2002] = -'sd58689;
    data[2003] =  'sd7344;
    data[2004] =  'sd19759;
    data[2005] =  'sd2452;
    data[2006] =  'sd61300;
    data[2007] =  'sd57931;
    data[2008] = -'sd26294;
    data[2009] = -'sd1986;
    data[2010] = -'sd49650;
    data[2011] =  'sd69478;
    data[2012] = -'sd65301;
    data[2013] =  'sd5885;
    data[2014] = -'sd16716;
    data[2015] =  'sd73623;
    data[2016] =  'sd38324;
    data[2017] = -'sd24946;
    data[2018] =  'sd31714;
    data[2019] = -'sd26355;
    data[2020] = -'sd3511;
    data[2021] =  'sd76066;
    data[2022] = -'sd64442;
    data[2023] =  'sd27360;
    data[2024] =  'sd28636;
    data[2025] =  'sd60536;
    data[2026] =  'sd38831;
    data[2027] = -'sd12271;
    data[2028] =  'sd20907;
    data[2029] =  'sd31152;
    data[2030] = -'sd40405;
    data[2031] = -'sd27079;
    data[2032] = -'sd21611;
    data[2033] = -'sd48752;
    data[2034] = -'sd71913;
    data[2035] =  'sd4426;
    data[2036] = -'sd53191;
    data[2037] = -'sd19047;
    data[2038] =  'sd15348;
    data[2039] =  'sd56018;
    data[2040] = -'sd74119;
    data[2041] = -'sd50724;
    data[2042] =  'sd42628;
    data[2043] = -'sd81187;
    data[2044] = -'sd63583;
    data[2045] =  'sd48835;
    data[2046] =  'sd73988;
    data[2047] =  'sd47449;
    data[2048] =  'sd39338;
    data[2049] =  'sd404;
    data[2050] =  'sd10100;
    data[2051] = -'sd75182;
    data[2052] = -'sd77299;
    data[2053] =  'sd33617;
    data[2054] =  'sd21220;
    data[2055] =  'sd38977;
    data[2056] = -'sd8621;
    data[2057] = -'sd51684;
    data[2058] =  'sd18628;
    data[2059] = -'sd25823;
    data[2060] =  'sd9789;
    data[2061] =  'sd80884;
    data[2062] =  'sd56008;
    data[2063] = -'sd74369;
    data[2064] = -'sd56974;
    data[2065] =  'sd50219;
    data[2066] = -'sd55253;
    data[2067] = -'sd70597;
    data[2068] =  'sd37326;
    data[2069] = -'sd49896;
    data[2070] =  'sd63328;
    data[2071] = -'sd55210;
    data[2072] = -'sd69522;
    data[2073] =  'sd64201;
    data[2074] = -'sd33385;
    data[2075] = -'sd15420;
    data[2076] = -'sd57818;
    data[2077] =  'sd29119;
    data[2078] =  'sd72611;
    data[2079] =  'sd13024;
    data[2080] = -'sd2082;
    data[2081] = -'sd52050;
    data[2082] =  'sd9478;
    data[2083] =  'sd73109;
    data[2084] =  'sd25474;
    data[2085] = -'sd18514;
    data[2086] =  'sd28673;
    data[2087] =  'sd61461;
    data[2088] =  'sd61956;
    data[2089] =  'sd74331;
    data[2090] =  'sd56024;
    data[2091] = -'sd73969;
    data[2092] = -'sd46974;
    data[2093] = -'sd27463;
    data[2094] = -'sd31211;
    data[2095] =  'sd38930;
    data[2096] = -'sd9796;
    data[2097] = -'sd81059;
    data[2098] = -'sd60383;
    data[2099] = -'sd35006;
    data[2100] = -'sd55945;
    data[2101] =  'sd75944;
    data[2102] = -'sd67492;
    data[2103] = -'sd48890;
    data[2104] = -'sd75363;
    data[2105] = -'sd81824;
    data[2106] = -'sd79508;
    data[2107] = -'sd21608;
    data[2108] = -'sd48677;
    data[2109] = -'sd70038;
    data[2110] =  'sd51301;
    data[2111] = -'sd28203;
    data[2112] = -'sd49711;
    data[2113] =  'sd67953;
    data[2114] =  'sd60415;
    data[2115] =  'sd35806;
    data[2116] =  'sd75945;
    data[2117] = -'sd67467;
    data[2118] = -'sd48265;
    data[2119] = -'sd59738;
    data[2120] = -'sd18881;
    data[2121] =  'sd19498;
    data[2122] = -'sd4073;
    data[2123] =  'sd62016;
    data[2124] =  'sd75831;
    data[2125] = -'sd70317;
    data[2126] =  'sd44326;
    data[2127] = -'sd38737;
    data[2128] =  'sd14621;
    data[2129] =  'sd37843;
    data[2130] = -'sd36971;
    data[2131] =  'sd58771;
    data[2132] = -'sd5294;
    data[2133] =  'sd31491;
    data[2134] = -'sd31930;
    data[2135] =  'sd20955;
    data[2136] =  'sd32352;
    data[2137] = -'sd10405;
    data[2138] =  'sd67557;
    data[2139] =  'sd50515;
    data[2140] = -'sd47853;
    data[2141] = -'sd49438;
    data[2142] =  'sd74778;
    data[2143] =  'sd67199;
    data[2144] =  'sd41565;
    data[2145] =  'sd56079;
    data[2146] = -'sd72594;
    data[2147] = -'sd12599;
    data[2148] =  'sd12707;
    data[2149] = -'sd10007;
    data[2150] =  'sd77507;
    data[2151] = -'sd28417;
    data[2152] = -'sd55061;
    data[2153] = -'sd65797;
    data[2154] = -'sd6515;
    data[2155] =  'sd966;
    data[2156] =  'sd24150;
    data[2157] = -'sd51614;
    data[2158] =  'sd20378;
    data[2159] =  'sd17927;
    data[2160] = -'sd43348;
    data[2161] =  'sd63187;
    data[2162] = -'sd58735;
    data[2163] =  'sd6194;
    data[2164] = -'sd8991;
    data[2165] = -'sd60934;
    data[2166] = -'sd48781;
    data[2167] = -'sd72638;
    data[2168] = -'sd13699;
    data[2169] = -'sd14793;
    data[2170] = -'sd42143;
    data[2171] = -'sd70529;
    data[2172] =  'sd39026;
    data[2173] = -'sd7396;
    data[2174] = -'sd21059;
    data[2175] = -'sd34952;
    data[2176] = -'sd54595;
    data[2177] = -'sd54147;
    data[2178] = -'sd42947;
    data[2179] =  'sd73212;
    data[2180] =  'sd28049;
    data[2181] =  'sd45861;
    data[2182] = -'sd362;
    data[2183] = -'sd9050;
    data[2184] = -'sd62409;
    data[2185] =  'sd78185;
    data[2186] = -'sd11467;
    data[2187] =  'sd41007;
    data[2188] =  'sd42129;
    data[2189] =  'sd70179;
    data[2190] = -'sd47776;
    data[2191] = -'sd47513;
    data[2192] = -'sd40938;
    data[2193] = -'sd40404;
    data[2194] = -'sd27054;
    data[2195] = -'sd20986;
    data[2196] = -'sd33127;
    data[2197] = -'sd8970;
    data[2198] = -'sd60409;
    data[2199] = -'sd35656;
    data[2200] = -'sd72195;
    data[2201] = -'sd2624;
    data[2202] = -'sd65600;
    data[2203] = -'sd1590;
    data[2204] = -'sd39750;
    data[2205] = -'sd10704;
    data[2206] =  'sd60082;
    data[2207] =  'sd27481;
    data[2208] =  'sd31661;
    data[2209] = -'sd27680;
    data[2210] = -'sd36636;
    data[2211] =  'sd67146;
    data[2212] =  'sd40240;
    data[2213] =  'sd22954;
    data[2214] = -'sd81514;
    data[2215] = -'sd71758;
    data[2216] =  'sd8301;
    data[2217] =  'sd43684;
    data[2218] = -'sd54787;
    data[2219] = -'sd58947;
    data[2220] =  'sd894;
    data[2221] =  'sd22350;
    data[2222] =  'sd67227;
    data[2223] =  'sd42265;
    data[2224] =  'sd73579;
    data[2225] =  'sd37224;
    data[2226] = -'sd52446;
    data[2227] = -'sd422;
    data[2228] = -'sd10550;
    data[2229] =  'sd63932;
    data[2230] = -'sd40110;
    data[2231] = -'sd19704;
    data[2232] = -'sd1077;
    data[2233] = -'sd26925;
    data[2234] = -'sd17761;
    data[2235] =  'sd47498;
    data[2236] =  'sd40563;
    data[2237] =  'sd31029;
    data[2238] = -'sd43480;
    data[2239] =  'sd59887;
    data[2240] =  'sd22606;
    data[2241] =  'sd73627;
    data[2242] =  'sd38424;
    data[2243] = -'sd22446;
    data[2244] = -'sd69627;
    data[2245] =  'sd61576;
    data[2246] =  'sd64831;
    data[2247] = -'sd17635;
    data[2248] =  'sd50648;
    data[2249] = -'sd44528;
    data[2250] =  'sd33687;
    data[2251] =  'sd22970;
    data[2252] = -'sd81114;
    data[2253] = -'sd61758;
    data[2254] = -'sd69381;
    data[2255] =  'sd67726;
    data[2256] =  'sd54740;
    data[2257] =  'sd57772;
    data[2258] = -'sd30269;
    data[2259] =  'sd62480;
    data[2260] = -'sd76410;
    data[2261] =  'sd55842;
    data[2262] = -'sd78519;
    data[2263] =  'sd3117;
    data[2264] =  'sd77925;
    data[2265] = -'sd17967;
    data[2266] =  'sd42348;
    data[2267] =  'sd75654;
    data[2268] = -'sd74742;
    data[2269] = -'sd66299;
    data[2270] = -'sd19065;
    data[2271] =  'sd14898;
    data[2272] =  'sd44768;
    data[2273] = -'sd27687;
    data[2274] = -'sd36811;
    data[2275] =  'sd62771;
    data[2276] = -'sd69135;
    data[2277] =  'sd73876;
    data[2278] =  'sd44649;
    data[2279] = -'sd30662;
    data[2280] =  'sd52655;
    data[2281] =  'sd5647;
    data[2282] = -'sd22666;
    data[2283] = -'sd75127;
    data[2284] = -'sd75924;
    data[2285] =  'sd67992;
    data[2286] =  'sd61390;
    data[2287] =  'sd60181;
    data[2288] =  'sd29956;
    data[2289] = -'sd70305;
    data[2290] =  'sd44626;
    data[2291] = -'sd31237;
    data[2292] =  'sd38280;
    data[2293] = -'sd26046;
    data[2294] =  'sd4214;
    data[2295] = -'sd58491;
    data[2296] =  'sd12294;
    data[2297] = -'sd20332;
    data[2298] = -'sd16777;
    data[2299] =  'sd72098;
    data[2300] =  'sd199;
    data[2301] =  'sd4975;
    data[2302] = -'sd39466;
    data[2303] = -'sd3604;
    data[2304] =  'sd73741;
    data[2305] =  'sd41274;
    data[2306] =  'sd48804;
    data[2307] =  'sd73213;
    data[2308] =  'sd28074;
    data[2309] =  'sd46486;
    data[2310] =  'sd15263;
    data[2311] =  'sd53893;
    data[2312] =  'sd36597;
    data[2313] = -'sd68121;
    data[2314] = -'sd64615;
    data[2315] =  'sd23035;
    data[2316] = -'sd79489;
    data[2317] = -'sd21133;
    data[2318] = -'sd36802;
    data[2319] =  'sd62996;
    data[2320] = -'sd63510;
    data[2321] =  'sd50660;
    data[2322] = -'sd44228;
    data[2323] =  'sd41187;
    data[2324] =  'sd46629;
    data[2325] =  'sd18838;
    data[2326] = -'sd20573;
    data[2327] = -'sd22802;
    data[2328] = -'sd78527;
    data[2329] =  'sd2917;
    data[2330] =  'sd72925;
    data[2331] =  'sd20874;
    data[2332] =  'sd30327;
    data[2333] = -'sd61030;
    data[2334] = -'sd51181;
    data[2335] =  'sd31203;
    data[2336] = -'sd39130;
    data[2337] =  'sd4796;
    data[2338] = -'sd43941;
    data[2339] =  'sd48362;
    data[2340] =  'sd62163;
    data[2341] =  'sd79506;
    data[2342] =  'sd21558;
    data[2343] =  'sd47427;
    data[2344] =  'sd38788;
    data[2345] = -'sd13346;
    data[2346] = -'sd5968;
    data[2347] =  'sd14641;
    data[2348] =  'sd38343;
    data[2349] = -'sd24471;
    data[2350] =  'sd43589;
    data[2351] = -'sd57162;
    data[2352] =  'sd45519;
    data[2353] = -'sd8912;
    data[2354] = -'sd58959;
    data[2355] =  'sd594;
    data[2356] =  'sd14850;
    data[2357] =  'sd43568;
    data[2358] = -'sd57687;
    data[2359] =  'sd32394;
    data[2360] = -'sd9355;
    data[2361] = -'sd70034;
    data[2362] =  'sd51401;
    data[2363] = -'sd25703;
    data[2364] =  'sd12789;
    data[2365] = -'sd7957;
    data[2366] = -'sd35084;
    data[2367] = -'sd57895;
    data[2368] =  'sd27194;
    data[2369] =  'sd24486;
    data[2370] = -'sd43214;
    data[2371] =  'sd66537;
    data[2372] =  'sd25015;
    data[2373] = -'sd29989;
    data[2374] =  'sd69480;
    data[2375] = -'sd65251;
    data[2376] =  'sd7135;
    data[2377] =  'sd14534;
    data[2378] =  'sd35668;
    data[2379] =  'sd72495;
    data[2380] =  'sd10124;
    data[2381] = -'sd74582;
    data[2382] = -'sd62299;
    data[2383] =  'sd80935;
    data[2384] =  'sd57283;
    data[2385] = -'sd42494;
    data[2386] = -'sd79304;
    data[2387] = -'sd16508;
    data[2388] =  'sd78823;
    data[2389] =  'sd4483;
    data[2390] = -'sd51766;
    data[2391] =  'sd16578;
    data[2392] = -'sd77073;
    data[2393] =  'sd39267;
    data[2394] = -'sd1371;
    data[2395] = -'sd34275;
    data[2396] = -'sd37670;
    data[2397] =  'sd41296;
    data[2398] =  'sd49354;
    data[2399] = -'sd76878;
    data[2400] =  'sd44142;
    data[2401] = -'sd43337;
    data[2402] =  'sd63462;
    data[2403] = -'sd51860;
    data[2404] =  'sd14228;
    data[2405] =  'sd28018;
    data[2406] =  'sd45086;
    data[2407] = -'sd19737;
    data[2408] = -'sd1902;
    data[2409] = -'sd47550;
    data[2410] = -'sd41863;
    data[2411] = -'sd63529;
    data[2412] =  'sd50185;
    data[2413] = -'sd56103;
    data[2414] =  'sd71994;
    data[2415] = -'sd2401;
    data[2416] = -'sd60025;
    data[2417] = -'sd26056;
    data[2418] =  'sd3964;
    data[2419] = -'sd64741;
    data[2420] =  'sd19885;
    data[2421] =  'sd5602;
    data[2422] = -'sd23791;
    data[2423] =  'sd60589;
    data[2424] =  'sd40156;
    data[2425] =  'sd20854;
    data[2426] =  'sd29827;
    data[2427] = -'sd73530;
    data[2428] = -'sd35999;
    data[2429] = -'sd80770;
    data[2430] = -'sd53158;
    data[2431] = -'sd18222;
    data[2432] =  'sd35973;
    data[2433] =  'sd80120;
    data[2434] =  'sd36908;
    data[2435] = -'sd60346;
    data[2436] = -'sd34081;
    data[2437] = -'sd32820;
    data[2438] = -'sd1295;
    data[2439] = -'sd32375;
    data[2440] =  'sd9830;
    data[2441] =  'sd81909;
    data[2442] =  'sd81633;
    data[2443] =  'sd74733;
    data[2444] =  'sd66074;
    data[2445] =  'sd13440;
    data[2446] =  'sd8318;
    data[2447] =  'sd44109;
    data[2448] = -'sd44162;
    data[2449] =  'sd42837;
    data[2450] = -'sd75962;
    data[2451] =  'sd67042;
    data[2452] =  'sd37640;
    data[2453] = -'sd42046;
    data[2454] = -'sd68104;
    data[2455] = -'sd64190;
    data[2456] =  'sd33660;
    data[2457] =  'sd22295;
    data[2458] =  'sd65852;
    data[2459] =  'sd7890;
    data[2460] =  'sd33409;
    data[2461] =  'sd16020;
    data[2462] =  'sd72818;
    data[2463] =  'sd18199;
    data[2464] = -'sd36548;
    data[2465] =  'sd69346;
    data[2466] = -'sd68601;
    data[2467] = -'sd76615;
    data[2468] =  'sd50717;
    data[2469] = -'sd42803;
    data[2470] =  'sd76812;
    data[2471] = -'sd45792;
    data[2472] =  'sd2087;
    data[2473] =  'sd52175;
    data[2474] = -'sd6353;
    data[2475] =  'sd5016;
    data[2476] = -'sd38441;
    data[2477] =  'sd22021;
    data[2478] =  'sd59002;
    data[2479] =  'sd481;
    data[2480] =  'sd12025;
    data[2481] = -'sd27057;
    data[2482] = -'sd21061;
    data[2483] = -'sd35002;
    data[2484] = -'sd55845;
    data[2485] =  'sd78444;
    data[2486] = -'sd4992;
    data[2487] =  'sd39041;
    data[2488] = -'sd7021;
    data[2489] = -'sd11684;
    data[2490] =  'sd35582;
    data[2491] =  'sd70345;
    data[2492] = -'sd43626;
    data[2493] =  'sd56237;
    data[2494] = -'sd68644;
    data[2495] = -'sd77690;
    data[2496] =  'sd23842;
    data[2497] = -'sd59314;
    data[2498] = -'sd8281;
    data[2499] = -'sd43184;
    data[2500] =  'sd67287;
    data[2501] =  'sd43765;
    data[2502] = -'sd52762;
    data[2503] = -'sd8322;
    data[2504] = -'sd44209;
    data[2505] =  'sd41662;
    data[2506] =  'sd58504;
    data[2507] = -'sd11969;
    data[2508] =  'sd28457;
    data[2509] =  'sd56061;
    data[2510] = -'sd73044;
    data[2511] = -'sd23849;
    data[2512] =  'sd59139;
    data[2513] =  'sd3906;
    data[2514] = -'sd66191;
    data[2515] = -'sd16365;
    data[2516] = -'sd81443;
    data[2517] = -'sd69983;
    data[2518] =  'sd52676;
    data[2519] =  'sd6172;
    data[2520] = -'sd9541;
    data[2521] = -'sd74684;
    data[2522] = -'sd64849;
    data[2523] =  'sd17185;
    data[2524] = -'sd61898;
    data[2525] = -'sd72881;
    data[2526] = -'sd19774;
    data[2527] = -'sd2827;
    data[2528] = -'sd70675;
    data[2529] =  'sd35376;
    data[2530] =  'sd65195;
    data[2531] = -'sd8535;
    data[2532] = -'sd49534;
    data[2533] =  'sd72378;
    data[2534] =  'sd7199;
    data[2535] =  'sd16134;
    data[2536] =  'sd75668;
    data[2537] = -'sd74392;
    data[2538] = -'sd57549;
    data[2539] =  'sd35844;
    data[2540] =  'sd76895;
    data[2541] = -'sd43717;
    data[2542] =  'sd53962;
    data[2543] =  'sd38322;
    data[2544] = -'sd24996;
    data[2545] =  'sd30464;
    data[2546] = -'sd57605;
    data[2547] =  'sd34444;
    data[2548] =  'sd41895;
    data[2549] =  'sd64329;
    data[2550] = -'sd30185;
    data[2551] =  'sd64580;
    data[2552] = -'sd23910;
    data[2553] =  'sd57614;
    data[2554] = -'sd34219;
    data[2555] = -'sd36270;
    data[2556] =  'sd76296;
    data[2557] = -'sd58692;
    data[2558] =  'sd7269;
    data[2559] =  'sd17884;
    data[2560] = -'sd44423;
    data[2561] =  'sd36312;
    data[2562] = -'sd75246;
    data[2563] = -'sd78899;
    data[2564] = -'sd6383;
    data[2565] =  'sd4266;
    data[2566] = -'sd57191;
    data[2567] =  'sd44794;
    data[2568] = -'sd27037;
    data[2569] = -'sd20561;
    data[2570] = -'sd22502;
    data[2571] = -'sd71027;
    data[2572] =  'sd26576;
    data[2573] =  'sd9036;
    data[2574] =  'sd62059;
    data[2575] =  'sd76906;
    data[2576] = -'sd43442;
    data[2577] =  'sd60837;
    data[2578] =  'sd46356;
    data[2579] =  'sd12013;
    data[2580] = -'sd27357;
    data[2581] = -'sd28561;
    data[2582] = -'sd58661;
    data[2583] =  'sd8044;
    data[2584] =  'sd37259;
    data[2585] = -'sd51571;
    data[2586] =  'sd21453;
    data[2587] =  'sd44802;
    data[2588] = -'sd26837;
    data[2589] = -'sd15561;
    data[2590] = -'sd61343;
    data[2591] = -'sd59006;
    data[2592] = -'sd581;
    data[2593] = -'sd14525;
    data[2594] = -'sd35443;
    data[2595] = -'sd66870;
    data[2596] = -'sd33340;
    data[2597] = -'sd14295;
    data[2598] = -'sd29693;
    data[2599] =  'sd76880;
    data[2600] = -'sd44092;
    data[2601] =  'sd44587;
    data[2602] = -'sd32212;
    data[2603] =  'sd13905;
    data[2604] =  'sd19943;
    data[2605] =  'sd7052;
    data[2606] =  'sd12459;
    data[2607] = -'sd16207;
    data[2608] = -'sd77493;
    data[2609] =  'sd28767;
    data[2610] =  'sd63811;
    data[2611] = -'sd43135;
    data[2612] =  'sd68512;
    data[2613] =  'sd74390;
    data[2614] =  'sd57499;
    data[2615] = -'sd37094;
    data[2616] =  'sd55696;
    data[2617] =  'sd81672;
    data[2618] =  'sd75708;
    data[2619] = -'sd73392;
    data[2620] = -'sd32549;
    data[2621] =  'sd5480;
    data[2622] = -'sd26841;
    data[2623] = -'sd15661;
    data[2624] = -'sd63843;
    data[2625] =  'sd42335;
    data[2626] =  'sd75329;
    data[2627] =  'sd80974;
    data[2628] =  'sd58258;
    data[2629] = -'sd18119;
    data[2630] =  'sd38548;
    data[2631] = -'sd19346;
    data[2632] =  'sd7873;
    data[2633] =  'sd32984;
    data[2634] =  'sd5395;
    data[2635] = -'sd28966;
    data[2636] = -'sd68786;
    data[2637] = -'sd81240;
    data[2638] = -'sd64908;
    data[2639] =  'sd15710;
    data[2640] =  'sd65068;
    data[2641] = -'sd11710;
    data[2642] =  'sd34932;
    data[2643] =  'sd54095;
    data[2644] =  'sd41647;
    data[2645] =  'sd58129;
    data[2646] = -'sd21344;
    data[2647] = -'sd42077;
    data[2648] = -'sd68879;
    data[2649] =  'sd80276;
    data[2650] =  'sd40808;
    data[2651] =  'sd37154;
    data[2652] = -'sd54196;
    data[2653] = -'sd44172;
    data[2654] =  'sd42587;
    data[2655] =  'sd81629;
    data[2656] =  'sd74633;
    data[2657] =  'sd63574;
    data[2658] = -'sd49060;
    data[2659] = -'sd79613;
    data[2660] = -'sd24233;
    data[2661] =  'sd49539;
    data[2662] = -'sd72253;
    data[2663] = -'sd4074;
    data[2664] =  'sd61991;
    data[2665] =  'sd75206;
    data[2666] =  'sd77899;
    data[2667] = -'sd18617;
    data[2668] =  'sd26098;
    data[2669] = -'sd2914;
    data[2670] = -'sd72850;
    data[2671] = -'sd18999;
    data[2672] =  'sd16548;
    data[2673] = -'sd77823;
    data[2674] =  'sd20517;
    data[2675] =  'sd21402;
    data[2676] =  'sd43527;
    data[2677] = -'sd58712;
    data[2678] =  'sd6769;
    data[2679] =  'sd5384;
    data[2680] = -'sd29241;
    data[2681] = -'sd75661;
    data[2682] =  'sd74567;
    data[2683] =  'sd61924;
    data[2684] =  'sd73531;
    data[2685] =  'sd36024;
    data[2686] =  'sd81395;
    data[2687] =  'sd68783;
    data[2688] =  'sd81165;
    data[2689] =  'sd63033;
    data[2690] = -'sd62585;
    data[2691] =  'sd73785;
    data[2692] =  'sd42374;
    data[2693] =  'sd76304;
    data[2694] = -'sd58492;
    data[2695] =  'sd12269;
    data[2696] = -'sd20957;
    data[2697] = -'sd32402;
    data[2698] =  'sd9155;
    data[2699] =  'sd65034;
    data[2700] = -'sd12560;
    data[2701] =  'sd13682;
    data[2702] =  'sd14368;
    data[2703] =  'sd31518;
    data[2704] = -'sd31255;
    data[2705] =  'sd37830;
    data[2706] = -'sd37296;
    data[2707] =  'sd50646;
    data[2708] = -'sd44578;
    data[2709] =  'sd32437;
    data[2710] = -'sd8280;
    data[2711] = -'sd43159;
    data[2712] =  'sd67912;
    data[2713] =  'sd59390;
    data[2714] =  'sd10181;
    data[2715] = -'sd73157;
    data[2716] = -'sd26674;
    data[2717] = -'sd11486;
    data[2718] =  'sd40532;
    data[2719] =  'sd30254;
    data[2720] = -'sd62855;
    data[2721] =  'sd67035;
    data[2722] =  'sd37465;
    data[2723] = -'sd46421;
    data[2724] = -'sd13638;
    data[2725] = -'sd13268;
    data[2726] = -'sd4018;
    data[2727] =  'sd63391;
    data[2728] = -'sd53635;
    data[2729] = -'sd30147;
    data[2730] =  'sd65530;
    data[2731] = -'sd160;
    data[2732] = -'sd4000;
    data[2733] =  'sd63841;
    data[2734] = -'sd42385;
    data[2735] = -'sd76579;
    data[2736] =  'sd51617;
    data[2737] = -'sd20303;
    data[2738] = -'sd16052;
    data[2739] = -'sd73618;
    data[2740] = -'sd38199;
    data[2741] =  'sd28071;
    data[2742] =  'sd46411;
    data[2743] =  'sd13388;
    data[2744] =  'sd7018;
    data[2745] =  'sd11609;
    data[2746] = -'sd37457;
    data[2747] =  'sd46621;
    data[2748] =  'sd18638;
    data[2749] = -'sd25573;
    data[2750] =  'sd16039;
    data[2751] =  'sd73293;
    data[2752] =  'sd30074;
    data[2753] = -'sd67355;
    data[2754] = -'sd45465;
    data[2755] =  'sd10262;
    data[2756] = -'sd71132;
    data[2757] =  'sd23951;
    data[2758] = -'sd56589;
    data[2759] =  'sd59844;
    data[2760] =  'sd21531;
    data[2761] =  'sd46752;
    data[2762] =  'sd21913;
    data[2763] =  'sd56302;
    data[2764] = -'sd67019;
    data[2765] = -'sd37065;
    data[2766] =  'sd56421;
    data[2767] = -'sd64044;
    data[2768] =  'sd37310;
    data[2769] = -'sd50296;
    data[2770] =  'sd53328;
    data[2771] =  'sd22472;
    data[2772] =  'sd70277;
    data[2773] = -'sd45326;
    data[2774] =  'sd13737;
    data[2775] =  'sd15743;
    data[2776] =  'sd65893;
    data[2777] =  'sd8915;
    data[2778] =  'sd59034;
    data[2779] =  'sd1281;
    data[2780] =  'sd32025;
    data[2781] = -'sd18580;
    data[2782] =  'sd27023;
    data[2783] =  'sd20211;
    data[2784] =  'sd13752;
    data[2785] =  'sd16118;
    data[2786] =  'sd75268;
    data[2787] =  'sd79449;
    data[2788] =  'sd20133;
    data[2789] =  'sd11802;
    data[2790] = -'sd32632;
    data[2791] =  'sd3405;
    data[2792] = -'sd78716;
    data[2793] = -'sd1808;
    data[2794] = -'sd45200;
    data[2795] =  'sd16887;
    data[2796] = -'sd69348;
    data[2797] =  'sd68551;
    data[2798] =  'sd75365;
    data[2799] =  'sd81874;
    data[2800] =  'sd80758;
    data[2801] =  'sd52858;
    data[2802] =  'sd10722;
    data[2803] = -'sd59632;
    data[2804] = -'sd16231;
    data[2805] = -'sd78093;
    data[2806] =  'sd13767;
    data[2807] =  'sd16493;
    data[2808] = -'sd79198;
    data[2809] = -'sd13858;
    data[2810] = -'sd18768;
    data[2811] =  'sd22323;
    data[2812] =  'sd66552;
    data[2813] =  'sd25390;
    data[2814] = -'sd20614;
    data[2815] = -'sd23827;
    data[2816] =  'sd59689;
    data[2817] =  'sd17656;
    data[2818] = -'sd50123;
    data[2819] =  'sd57653;
    data[2820] = -'sd33244;
    data[2821] = -'sd11895;
    data[2822] =  'sd30307;
    data[2823] = -'sd61530;
    data[2824] = -'sd63681;
    data[2825] =  'sd46385;
    data[2826] =  'sd12738;
    data[2827] = -'sd9232;
    data[2828] = -'sd66959;
    data[2829] = -'sd35565;
    data[2830] = -'sd69920;
    data[2831] =  'sd54251;
    data[2832] =  'sd45547;
    data[2833] = -'sd8212;
    data[2834] = -'sd41459;
    data[2835] = -'sd53429;
    data[2836] = -'sd24997;
    data[2837] =  'sd30439;
    data[2838] = -'sd58230;
    data[2839] =  'sd18819;
    data[2840] = -'sd21048;
    data[2841] = -'sd34677;
    data[2842] = -'sd47720;
    data[2843] = -'sd46113;
    data[2844] = -'sd5938;
    data[2845] =  'sd15391;
    data[2846] =  'sd57093;
    data[2847] = -'sd47244;
    data[2848] = -'sd34213;
    data[2849] = -'sd36120;
    data[2850] =  'sd80046;
    data[2851] =  'sd35058;
    data[2852] =  'sd57245;
    data[2853] = -'sd43444;
    data[2854] =  'sd60787;
    data[2855] =  'sd45106;
    data[2856] = -'sd19237;
    data[2857] =  'sd10598;
    data[2858] = -'sd62732;
    data[2859] =  'sd70110;
    data[2860] = -'sd49501;
    data[2861] =  'sd73203;
    data[2862] =  'sd27824;
    data[2863] =  'sd40236;
    data[2864] =  'sd22854;
    data[2865] =  'sd79827;
    data[2866] =  'sd29583;
    data[2867] = -'sd79630;
    data[2868] = -'sd24658;
    data[2869] =  'sd38914;
    data[2870] = -'sd10196;
    data[2871] =  'sd72782;
    data[2872] =  'sd17299;
    data[2873] = -'sd59048;
    data[2874] = -'sd1631;
    data[2875] = -'sd40775;
    data[2876] = -'sd36329;
    data[2877] =  'sd74821;
    data[2878] =  'sd68274;
    data[2879] =  'sd68440;
    data[2880] =  'sd72590;
    data[2881] =  'sd12499;
    data[2882] = -'sd15207;
    data[2883] = -'sd52493;
    data[2884] = -'sd1597;
    data[2885] = -'sd39925;
    data[2886] = -'sd15079;
    data[2887] = -'sd49293;
    data[2888] =  'sd78403;
    data[2889] = -'sd6017;
    data[2890] =  'sd13416;
    data[2891] =  'sd7718;
    data[2892] =  'sd29109;
    data[2893] =  'sd72361;
    data[2894] =  'sd6774;
    data[2895] =  'sd5509;
    data[2896] = -'sd26116;
    data[2897] =  'sd2464;
    data[2898] =  'sd61600;
    data[2899] =  'sd65431;
    data[2900] = -'sd2635;
    data[2901] = -'sd65875;
    data[2902] = -'sd8465;
    data[2903] = -'sd47784;
    data[2904] = -'sd47713;
    data[2905] = -'sd45938;
    data[2906] = -'sd1563;
    data[2907] = -'sd39075;
    data[2908] =  'sd6171;
    data[2909] = -'sd9566;
    data[2910] = -'sd75309;
    data[2911] = -'sd80474;
    data[2912] = -'sd45758;
    data[2913] =  'sd2937;
    data[2914] =  'sd73425;
    data[2915] =  'sd33374;
    data[2916] =  'sd15145;
    data[2917] =  'sd50943;
    data[2918] = -'sd37153;
    data[2919] =  'sd54221;
    data[2920] =  'sd44797;
    data[2921] = -'sd26962;
    data[2922] = -'sd18686;
    data[2923] =  'sd24373;
    data[2924] = -'sd46039;
    data[2925] = -'sd4088;
    data[2926] =  'sd61641;
    data[2927] =  'sd66456;
    data[2928] =  'sd22990;
    data[2929] = -'sd80614;
    data[2930] = -'sd49258;
    data[2931] =  'sd79278;
    data[2932] =  'sd15858;
    data[2933] =  'sd68768;
    data[2934] =  'sd80790;
    data[2935] =  'sd53658;
    data[2936] =  'sd30722;
    data[2937] = -'sd51155;
    data[2938] =  'sd31853;
    data[2939] = -'sd22880;
    data[2940] = -'sd80477;
    data[2941] = -'sd45833;
    data[2942] =  'sd1062;
    data[2943] =  'sd26550;
    data[2944] =  'sd8386;
    data[2945] =  'sd45809;
    data[2946] = -'sd1662;
    data[2947] = -'sd41550;
    data[2948] = -'sd55704;
    data[2949] = -'sd81872;
    data[2950] = -'sd80708;
    data[2951] = -'sd51608;
    data[2952] =  'sd20528;
    data[2953] =  'sd21677;
    data[2954] =  'sd50402;
    data[2955] = -'sd50678;
    data[2956] =  'sd43778;
    data[2957] = -'sd52437;
    data[2958] = -'sd197;
    data[2959] = -'sd4925;
    data[2960] =  'sd40716;
    data[2961] =  'sd34854;
    data[2962] =  'sd52145;
    data[2963] = -'sd7103;
    data[2964] = -'sd13734;
    data[2965] = -'sd15668;
    data[2966] = -'sd64018;
    data[2967] =  'sd37960;
    data[2968] = -'sd34046;
    data[2969] = -'sd31945;
    data[2970] =  'sd20580;
    data[2971] =  'sd22977;
    data[2972] = -'sd80939;
    data[2973] = -'sd57383;
    data[2974] =  'sd39994;
    data[2975] =  'sd16804;
    data[2976] = -'sd71423;
    data[2977] =  'sd16676;
    data[2978] = -'sd74623;
    data[2979] = -'sd63324;
    data[2980] =  'sd55310;
    data[2981] =  'sd72022;
    data[2982] = -'sd1701;
    data[2983] = -'sd42525;
    data[2984] = -'sd80079;
    data[2985] = -'sd35883;
    data[2986] = -'sd77870;
    data[2987] =  'sd19342;
    data[2988] = -'sd7973;
    data[2989] = -'sd35484;
    data[2990] = -'sd67895;
    data[2991] = -'sd58965;
    data[2992] =  'sd444;
    data[2993] =  'sd11100;
    data[2994] = -'sd50182;
    data[2995] =  'sd56178;
    data[2996] = -'sd70119;
    data[2997] =  'sd49276;
    data[2998] = -'sd78828;
    data[2999] = -'sd4608;
    data[3000] =  'sd48641;
    data[3001] =  'sd69138;
    data[3002] = -'sd73801;
    data[3003] = -'sd42774;
    data[3004] =  'sd77537;
    data[3005] = -'sd27667;
    data[3006] = -'sd36311;
    data[3007] =  'sd75271;
    data[3008] =  'sd79524;
    data[3009] =  'sd22008;
    data[3010] =  'sd58677;
    data[3011] = -'sd7644;
    data[3012] = -'sd27259;
    data[3013] = -'sd26111;
    data[3014] =  'sd2589;
    data[3015] =  'sd64725;
    data[3016] = -'sd20285;
    data[3017] = -'sd15602;
    data[3018] = -'sd62368;
    data[3019] =  'sd79210;
    data[3020] =  'sd14158;
    data[3021] =  'sd26268;
    data[3022] =  'sd1336;
    data[3023] =  'sd33400;
    data[3024] =  'sd15795;
    data[3025] =  'sd67193;
    data[3026] =  'sd41415;
    data[3027] =  'sd52329;
    data[3028] = -'sd2503;
    data[3029] = -'sd62575;
    data[3030] =  'sd74035;
    data[3031] =  'sd48624;
    data[3032] =  'sd68713;
    data[3033] =  'sd79415;
    data[3034] =  'sd19283;
    data[3035] = -'sd9448;
    data[3036] = -'sd72359;
    data[3037] = -'sd6724;
    data[3038] = -'sd4259;
    data[3039] =  'sd57366;
    data[3040] = -'sd40419;
    data[3041] = -'sd27429;
    data[3042] = -'sd30361;
    data[3043] =  'sd60180;
    data[3044] =  'sd29931;
    data[3045] = -'sd70930;
    data[3046] =  'sd29001;
    data[3047] =  'sd69661;
    data[3048] = -'sd60726;
    data[3049] = -'sd43581;
    data[3050] =  'sd57362;
    data[3051] = -'sd40519;
    data[3052] = -'sd29929;
    data[3053] =  'sd70980;
    data[3054] = -'sd27751;
    data[3055] = -'sd38411;
    data[3056] =  'sd22771;
    data[3057] =  'sd77752;
    data[3058] = -'sd22292;
    data[3059] = -'sd65777;
    data[3060] = -'sd6015;
    data[3061] =  'sd13466;
    data[3062] =  'sd8968;
    data[3063] =  'sd60359;
    data[3064] =  'sd34406;
    data[3065] =  'sd40945;
    data[3066] =  'sd40579;
    data[3067] =  'sd31429;
    data[3068] = -'sd33480;
    data[3069] = -'sd17795;
    data[3070] =  'sd46648;
    data[3071] =  'sd19313;
    data[3072] = -'sd8698;
    data[3073] = -'sd53609;
    data[3074] = -'sd29497;
    data[3075] =  'sd81780;
    data[3076] =  'sd78408;
    data[3077] = -'sd5892;
    data[3078] =  'sd16541;
    data[3079] = -'sd77998;
    data[3080] =  'sd16142;
    data[3081] =  'sd75868;
    data[3082] = -'sd69392;
    data[3083] =  'sd67451;
    data[3084] =  'sd47865;
    data[3085] =  'sd49738;
    data[3086] = -'sd67278;
    data[3087] = -'sd43540;
    data[3088] =  'sd58387;
    data[3089] = -'sd14894;
    data[3090] = -'sd44668;
    data[3091] =  'sd30187;
    data[3092] = -'sd64530;
    data[3093] =  'sd25160;
    data[3094] = -'sd26364;
    data[3095] = -'sd3736;
    data[3096] =  'sd70441;
    data[3097] = -'sd41226;
    data[3098] = -'sd47604;
    data[3099] = -'sd43213;
    data[3100] =  'sd66562;
    data[3101] =  'sd25640;
    data[3102] = -'sd14364;
    data[3103] = -'sd31418;
    data[3104] =  'sd33755;
    data[3105] =  'sd24670;
    data[3106] = -'sd38614;
    data[3107] =  'sd17696;
    data[3108] = -'sd49123;
    data[3109] = -'sd81188;
    data[3110] = -'sd63608;
    data[3111] =  'sd48210;
    data[3112] =  'sd58363;
    data[3113] = -'sd15494;
    data[3114] = -'sd59668;
    data[3115] = -'sd17131;
    data[3116] =  'sd63248;
    data[3117] = -'sd57210;
    data[3118] =  'sd44319;
    data[3119] = -'sd38912;
    data[3120] =  'sd10246;
    data[3121] = -'sd71532;
    data[3122] =  'sd13951;
    data[3123] =  'sd21093;
    data[3124] =  'sd35802;
    data[3125] =  'sd75845;
    data[3126] = -'sd69967;
    data[3127] =  'sd53076;
    data[3128] =  'sd16172;
    data[3129] =  'sd76618;
    data[3130] = -'sd50642;
    data[3131] =  'sd44678;
    data[3132] = -'sd29937;
    data[3133] =  'sd70780;
    data[3134] = -'sd32751;
    data[3135] =  'sd430;
    data[3136] =  'sd10750;
    data[3137] = -'sd58932;
    data[3138] =  'sd1269;
    data[3139] =  'sd31725;
    data[3140] = -'sd26080;
    data[3141] =  'sd3364;
    data[3142] = -'sd79741;
    data[3143] = -'sd27433;
    data[3144] = -'sd30461;
    data[3145] =  'sd57680;
    data[3146] = -'sd32569;
    data[3147] =  'sd4980;
    data[3148] = -'sd39341;
    data[3149] = -'sd479;
    data[3150] = -'sd11975;
    data[3151] =  'sd28307;
    data[3152] =  'sd52311;
    data[3153] = -'sd2953;
    data[3154] = -'sd73825;
    data[3155] = -'sd43374;
    data[3156] =  'sd62537;
    data[3157] = -'sd74985;
    data[3158] = -'sd72374;
    data[3159] = -'sd7099;
    data[3160] = -'sd13634;
    data[3161] = -'sd13168;
    data[3162] = -'sd1518;
    data[3163] = -'sd37950;
    data[3164] =  'sd34296;
    data[3165] =  'sd38195;
    data[3166] = -'sd28171;
    data[3167] = -'sd48911;
    data[3168] = -'sd75888;
    data[3169] =  'sd68892;
    data[3170] = -'sd79951;
    data[3171] = -'sd32683;
    data[3172] =  'sd2130;
    data[3173] =  'sd53250;
    data[3174] =  'sd20522;
    data[3175] =  'sd21527;
    data[3176] =  'sd46652;
    data[3177] =  'sd19413;
    data[3178] = -'sd6198;
    data[3179] =  'sd8891;
    data[3180] =  'sd58434;
    data[3181] = -'sd13719;
    data[3182] = -'sd15293;
    data[3183] = -'sd54643;
    data[3184] = -'sd55347;
    data[3185] = -'sd72947;
    data[3186] = -'sd21424;
    data[3187] = -'sd44077;
    data[3188] =  'sd44962;
    data[3189] = -'sd22837;
    data[3190] = -'sd79402;
    data[3191] = -'sd18958;
    data[3192] =  'sd17573;
    data[3193] = -'sd52198;
    data[3194] =  'sd5778;
    data[3195] = -'sd19391;
    data[3196] =  'sd6748;
    data[3197] =  'sd4859;
    data[3198] = -'sd42366;
    data[3199] = -'sd76104;
    data[3200] =  'sd63492;
    data[3201] = -'sd51110;
    data[3202] =  'sd32978;
    data[3203] =  'sd5245;
    data[3204] = -'sd32716;
    data[3205] =  'sd1305;
    data[3206] =  'sd32625;
    data[3207] = -'sd3580;
    data[3208] =  'sd74341;
    data[3209] =  'sd56274;
    data[3210] = -'sd67719;
    data[3211] = -'sd54565;
    data[3212] = -'sd53397;
    data[3213] = -'sd24197;
    data[3214] =  'sd50439;
    data[3215] = -'sd49753;
    data[3216] =  'sd66903;
    data[3217] =  'sd34165;
    data[3218] =  'sd34920;
    data[3219] =  'sd53795;
    data[3220] =  'sd34147;
    data[3221] =  'sd34470;
    data[3222] =  'sd42545;
    data[3223] =  'sd80579;
    data[3224] =  'sd48383;
    data[3225] =  'sd62688;
    data[3226] = -'sd71210;
    data[3227] =  'sd22001;
    data[3228] =  'sd58502;
    data[3229] = -'sd12019;
    data[3230] =  'sd27207;
    data[3231] =  'sd24811;
    data[3232] = -'sd35089;
    data[3233] = -'sd58020;
    data[3234] =  'sd24069;
    data[3235] = -'sd53639;
    data[3236] = -'sd30247;
    data[3237] =  'sd63030;
    data[3238] = -'sd62660;
    data[3239] =  'sd71910;
    data[3240] = -'sd4501;
    data[3241] =  'sd51316;
    data[3242] = -'sd27828;
    data[3243] = -'sd40336;
    data[3244] = -'sd25354;
    data[3245] =  'sd21514;
    data[3246] =  'sd46327;
    data[3247] =  'sd11288;
    data[3248] = -'sd45482;
    data[3249] =  'sd9837;
    data[3250] = -'sd81757;
    data[3251] = -'sd77833;
    data[3252] =  'sd20267;
    data[3253] =  'sd15152;
    data[3254] =  'sd51118;
    data[3255] = -'sd32778;
    data[3256] = -'sd245;
    data[3257] = -'sd6125;
    data[3258] =  'sd10716;
    data[3259] = -'sd59782;
    data[3260] = -'sd19981;
    data[3261] = -'sd8002;
    data[3262] = -'sd36209;
    data[3263] =  'sd77821;
    data[3264] = -'sd20567;
    data[3265] = -'sd22652;
    data[3266] = -'sd74777;
    data[3267] = -'sd67174;
    data[3268] = -'sd40940;
    data[3269] = -'sd40454;
    data[3270] = -'sd28304;
    data[3271] = -'sd52236;
    data[3272] =  'sd4828;
    data[3273] = -'sd43141;
    data[3274] =  'sd68362;
    data[3275] =  'sd70640;
    data[3276] = -'sd36251;
    data[3277] =  'sd76771;
    data[3278] = -'sd46817;
    data[3279] = -'sd23538;
    data[3280] =  'sd66914;
    data[3281] =  'sd34440;
    data[3282] =  'sd41795;
    data[3283] =  'sd61829;
    data[3284] =  'sd71156;
    data[3285] = -'sd23351;
    data[3286] =  'sd71589;
    data[3287] = -'sd12526;
    data[3288] =  'sd14532;
    data[3289] =  'sd35618;
    data[3290] =  'sd71245;
    data[3291] = -'sd21126;
    data[3292] = -'sd36627;
    data[3293] =  'sd67371;
    data[3294] =  'sd45865;
    data[3295] = -'sd262;
    data[3296] = -'sd6550;
    data[3297] =  'sd91;
    data[3298] =  'sd2275;
    data[3299] =  'sd56875;
    data[3300] = -'sd52694;
    data[3301] = -'sd6622;
    data[3302] = -'sd1709;
    data[3303] = -'sd42725;
    data[3304] =  'sd78762;
    data[3305] =  'sd2958;
    data[3306] =  'sd73950;
    data[3307] =  'sd46499;
    data[3308] =  'sd15588;
    data[3309] =  'sd62018;
    data[3310] =  'sd75881;
    data[3311] = -'sd69067;
    data[3312] =  'sd75576;
    data[3313] = -'sd76692;
    data[3314] =  'sd48792;
    data[3315] =  'sd72913;
    data[3316] =  'sd20574;
    data[3317] =  'sd22827;
    data[3318] =  'sd79152;
    data[3319] =  'sd12708;
    data[3320] = -'sd9982;
    data[3321] =  'sd78132;
    data[3322] = -'sd12792;
    data[3323] =  'sd7882;
    data[3324] =  'sd33209;
    data[3325] =  'sd11020;
    data[3326] = -'sd52182;
    data[3327] =  'sd6178;
    data[3328] = -'sd9391;
    data[3329] = -'sd70934;
    data[3330] =  'sd28901;
    data[3331] =  'sd67161;
    data[3332] =  'sd40615;
    data[3333] =  'sd32329;
    data[3334] = -'sd10980;
    data[3335] =  'sd53182;
    data[3336] =  'sd18822;
    data[3337] = -'sd20973;
    data[3338] = -'sd32802;
    data[3339] = -'sd845;
    data[3340] = -'sd21125;
    data[3341] = -'sd36602;
    data[3342] =  'sd67996;
    data[3343] =  'sd61490;
    data[3344] =  'sd62681;
    data[3345] = -'sd71385;
    data[3346] =  'sd17626;
    data[3347] = -'sd50873;
    data[3348] =  'sd38903;
    data[3349] = -'sd10471;
    data[3350] =  'sd65907;
    data[3351] =  'sd9265;
    data[3352] =  'sd67784;
    data[3353] =  'sd56190;
    data[3354] = -'sd69819;
    data[3355] =  'sd56776;
    data[3356] = -'sd55169;
    data[3357] = -'sd68497;
    data[3358] = -'sd74015;
    data[3359] = -'sd48124;
    data[3360] = -'sd56213;
    data[3361] =  'sd69244;
    data[3362] = -'sd71151;
    data[3363] =  'sd23476;
    data[3364] = -'sd68464;
    data[3365] = -'sd73190;
    data[3366] = -'sd27499;
    data[3367] = -'sd32111;
    data[3368] =  'sd16430;
    data[3369] = -'sd80773;
    data[3370] = -'sd53233;
    data[3371] = -'sd20097;
    data[3372] = -'sd10902;
    data[3373] =  'sd55132;
    data[3374] =  'sd67572;
    data[3375] =  'sd50890;
    data[3376] = -'sd38478;
    data[3377] =  'sd21096;
    data[3378] =  'sd35877;
    data[3379] =  'sd77720;
    data[3380] = -'sd23092;
    data[3381] =  'sd78064;
    data[3382] = -'sd14492;
    data[3383] = -'sd34618;
    data[3384] = -'sd46245;
    data[3385] = -'sd9238;
    data[3386] = -'sd67109;
    data[3387] = -'sd39315;
    data[3388] =  'sd171;
    data[3389] =  'sd4275;
    data[3390] = -'sd56966;
    data[3391] =  'sd50419;
    data[3392] = -'sd50253;
    data[3393] =  'sd54403;
    data[3394] =  'sd49347;
    data[3395] = -'sd77053;
    data[3396] =  'sd39767;
    data[3397] =  'sd11129;
    data[3398] = -'sd49457;
    data[3399] =  'sd74303;
    data[3400] =  'sd55324;
    data[3401] =  'sd72372;
    data[3402] =  'sd7049;
    data[3403] =  'sd12384;
    data[3404] = -'sd18082;
    data[3405] =  'sd39473;
    data[3406] =  'sd3779;
    data[3407] = -'sd69366;
    data[3408] =  'sd68101;
    data[3409] =  'sd64115;
    data[3410] = -'sd35535;
    data[3411] = -'sd69170;
    data[3412] =  'sd73001;
    data[3413] =  'sd22774;
    data[3414] =  'sd77827;
    data[3415] = -'sd20417;
    data[3416] = -'sd18902;
    data[3417] =  'sd18973;
    data[3418] = -'sd17198;
    data[3419] =  'sd61573;
    data[3420] =  'sd64756;
    data[3421] = -'sd19510;
    data[3422] =  'sd3773;
    data[3423] = -'sd69516;
    data[3424] =  'sd64351;
    data[3425] = -'sd29635;
    data[3426] =  'sd78330;
    data[3427] = -'sd7842;
    data[3428] = -'sd32209;
    data[3429] =  'sd13980;
    data[3430] =  'sd21818;
    data[3431] =  'sd53927;
    data[3432] =  'sd37447;
    data[3433] = -'sd46871;
    data[3434] = -'sd24888;
    data[3435] =  'sd33164;
    data[3436] =  'sd9895;
    data[3437] = -'sd80307;
    data[3438] = -'sd41583;
    data[3439] = -'sd56529;
    data[3440] =  'sd61344;
    data[3441] =  'sd59031;
    data[3442] =  'sd1206;
    data[3443] =  'sd30150;
    data[3444] = -'sd65455;
    data[3445] =  'sd2035;
    data[3446] =  'sd50875;
    data[3447] = -'sd38853;
    data[3448] =  'sd11721;
    data[3449] = -'sd34657;
    data[3450] = -'sd47220;
    data[3451] = -'sd33613;
    data[3452] = -'sd21120;
    data[3453] = -'sd36477;
    data[3454] =  'sd71121;
    data[3455] = -'sd24226;
    data[3456] =  'sd49714;
    data[3457] = -'sd67878;
    data[3458] = -'sd58540;
    data[3459] =  'sd11069;
    data[3460] = -'sd50957;
    data[3461] =  'sd36803;
    data[3462] = -'sd62971;
    data[3463] =  'sd64135;
    data[3464] = -'sd35035;
    data[3465] = -'sd56670;
    data[3466] =  'sd57819;
    data[3467] = -'sd29094;
    data[3468] = -'sd71986;
    data[3469] =  'sd2601;
    data[3470] =  'sd65025;
    data[3471] = -'sd12785;
    data[3472] =  'sd8057;
    data[3473] =  'sd37584;
    data[3474] = -'sd43446;
    data[3475] =  'sd60737;
    data[3476] =  'sd43856;
    data[3477] = -'sd50487;
    data[3478] =  'sd48553;
    data[3479] =  'sd66938;
    data[3480] =  'sd35040;
    data[3481] =  'sd56795;
    data[3482] = -'sd54694;
    data[3483] = -'sd56622;
    data[3484] =  'sd59019;
    data[3485] =  'sd906;
    data[3486] =  'sd22650;
    data[3487] =  'sd74727;
    data[3488] =  'sd65924;
    data[3489] =  'sd9690;
    data[3490] =  'sd78409;
    data[3491] = -'sd5867;
    data[3492] =  'sd17166;
    data[3493] = -'sd62373;
    data[3494] =  'sd79085;
    data[3495] =  'sd11033;
    data[3496] = -'sd51857;
    data[3497] =  'sd14303;
    data[3498] =  'sd29893;
    data[3499] = -'sd71880;
    data[3500] =  'sd5251;
    data[3501] = -'sd32566;
    data[3502] =  'sd5055;
    data[3503] = -'sd37466;
    data[3504] =  'sd46396;
    data[3505] =  'sd13013;
    data[3506] = -'sd2357;
    data[3507] = -'sd58925;
    data[3508] =  'sd1444;
    data[3509] =  'sd36100;
    data[3510] = -'sd80546;
    data[3511] = -'sd47558;
    data[3512] = -'sd42063;
    data[3513] = -'sd68529;
    data[3514] = -'sd74815;
    data[3515] = -'sd68124;
    data[3516] = -'sd64690;
    data[3517] =  'sd21160;
    data[3518] =  'sd37477;
    data[3519] = -'sd46121;
    data[3520] = -'sd6138;
    data[3521] =  'sd10391;
    data[3522] = -'sd67907;
    data[3523] = -'sd59265;
    data[3524] = -'sd7056;
    data[3525] = -'sd12559;
    data[3526] =  'sd13707;
    data[3527] =  'sd14993;
    data[3528] =  'sd47143;
    data[3529] =  'sd31688;
    data[3530] = -'sd27005;
    data[3531] = -'sd19761;
    data[3532] = -'sd2502;
    data[3533] = -'sd62550;
    data[3534] =  'sd74660;
    data[3535] =  'sd64249;
    data[3536] = -'sd32185;
    data[3537] =  'sd14580;
    data[3538] =  'sd36818;
    data[3539] = -'sd62596;
    data[3540] =  'sd73510;
    data[3541] =  'sd35499;
    data[3542] =  'sd68270;
    data[3543] =  'sd68340;
    data[3544] =  'sd70090;
    data[3545] = -'sd50001;
    data[3546] =  'sd60703;
    data[3547] =  'sd43006;
    data[3548] = -'sd71737;
    data[3549] =  'sd8826;
    data[3550] =  'sd56809;
    data[3551] = -'sd54344;
    data[3552] = -'sd47872;
    data[3553] = -'sd49913;
    data[3554] =  'sd62903;
    data[3555] = -'sd65835;
    data[3556] = -'sd7465;
    data[3557] = -'sd22784;
    data[3558] = -'sd78077;
    data[3559] =  'sd14167;
    data[3560] =  'sd26493;
    data[3561] =  'sd6961;
    data[3562] =  'sd10184;
    data[3563] = -'sd73082;
    data[3564] = -'sd24799;
    data[3565] =  'sd35389;
    data[3566] =  'sd65520;
    data[3567] = -'sd410;
    data[3568] = -'sd10250;
    data[3569] =  'sd71432;
    data[3570] = -'sd16451;
    data[3571] =  'sd80248;
    data[3572] =  'sd40108;
    data[3573] =  'sd19654;
    data[3574] = -'sd173;
    data[3575] = -'sd4325;
    data[3576] =  'sd55716;
    data[3577] = -'sd81669;
    data[3578] = -'sd75633;
    data[3579] =  'sd75267;
    data[3580] =  'sd79424;
    data[3581] =  'sd19508;
    data[3582] = -'sd3823;
    data[3583] =  'sd68266;
    data[3584] =  'sd68240;
    data[3585] =  'sd67590;
    data[3586] =  'sd51340;
    data[3587] = -'sd27228;
    data[3588] = -'sd25336;
    data[3589] =  'sd21964;
    data[3590] =  'sd57577;
    data[3591] = -'sd35144;
    data[3592] = -'sd59395;
    data[3593] = -'sd10306;
    data[3594] =  'sd70032;
    data[3595] = -'sd51451;
    data[3596] =  'sd24453;
    data[3597] = -'sd44039;
    data[3598] =  'sd45912;
    data[3599] =  'sd913;
    data[3600] =  'sd22825;
    data[3601] =  'sd79102;
    data[3602] =  'sd11458;
    data[3603] = -'sd41232;
    data[3604] = -'sd47754;
    data[3605] = -'sd46963;
    data[3606] = -'sd27188;
    data[3607] = -'sd24336;
    data[3608] =  'sd46964;
    data[3609] =  'sd27213;
    data[3610] =  'sd24961;
    data[3611] = -'sd31339;
    data[3612] =  'sd35730;
    data[3613] =  'sd74045;
    data[3614] =  'sd48874;
    data[3615] =  'sd74963;
    data[3616] =  'sd71824;
    data[3617] = -'sd6651;
    data[3618] = -'sd2434;
    data[3619] = -'sd60850;
    data[3620] = -'sd46681;
    data[3621] = -'sd20138;
    data[3622] = -'sd11927;
    data[3623] =  'sd29507;
    data[3624] = -'sd81530;
    data[3625] = -'sd72158;
    data[3626] = -'sd1699;
    data[3627] = -'sd42475;
    data[3628] = -'sd78829;
    data[3629] = -'sd4633;
    data[3630] =  'sd48016;
    data[3631] =  'sd53513;
    data[3632] =  'sd27097;
    data[3633] =  'sd22061;
    data[3634] =  'sd60002;
    data[3635] =  'sd25481;
    data[3636] = -'sd18339;
    data[3637] =  'sd33048;
    data[3638] =  'sd6995;
    data[3639] =  'sd11034;
    data[3640] = -'sd51832;
    data[3641] =  'sd14928;
    data[3642] =  'sd45518;
    data[3643] = -'sd8937;
    data[3644] = -'sd59584;
    data[3645] = -'sd15031;
    data[3646] = -'sd48093;
    data[3647] = -'sd55438;
    data[3648] = -'sd75222;
    data[3649] = -'sd78299;
    data[3650] =  'sd8617;
    data[3651] =  'sd51584;
    data[3652] = -'sd21128;
    data[3653] = -'sd36677;
    data[3654] =  'sd66121;
    data[3655] =  'sd14615;
    data[3656] =  'sd37693;
    data[3657] = -'sd40721;
    data[3658] = -'sd34979;
    data[3659] = -'sd55270;
    data[3660] = -'sd71022;
    data[3661] =  'sd26701;
    data[3662] =  'sd12161;
    data[3663] = -'sd23657;
    data[3664] =  'sd63939;
    data[3665] = -'sd39935;
    data[3666] = -'sd15329;
    data[3667] = -'sd55543;
    data[3668] = -'sd77847;
    data[3669] =  'sd19917;
    data[3670] =  'sd6402;
    data[3671] = -'sd3791;
    data[3672] =  'sd69066;
    data[3673] = -'sd75601;
    data[3674] =  'sd76067;
    data[3675] = -'sd64417;
    data[3676] =  'sd27985;
    data[3677] =  'sd44261;
    data[3678] = -'sd40362;
    data[3679] = -'sd26004;
    data[3680] =  'sd5264;
    data[3681] = -'sd32241;
    data[3682] =  'sd13180;
    data[3683] =  'sd1818;
    data[3684] =  'sd45450;
    data[3685] = -'sd10637;
    data[3686] =  'sd61757;
    data[3687] =  'sd69356;
    data[3688] = -'sd68351;
    data[3689] = -'sd70365;
    data[3690] =  'sd43126;
    data[3691] = -'sd68737;
    data[3692] = -'sd80015;
    data[3693] = -'sd34283;
    data[3694] = -'sd37870;
    data[3695] =  'sd36296;
    data[3696] = -'sd75646;
    data[3697] =  'sd74942;
    data[3698] =  'sd71299;
    data[3699] = -'sd19776;
    data[3700] = -'sd2877;
    data[3701] = -'sd71925;
    data[3702] =  'sd4126;
    data[3703] = -'sd60691;
    data[3704] = -'sd42706;
    data[3705] =  'sd79237;
    data[3706] =  'sd14833;
    data[3707] =  'sd43143;
    data[3708] = -'sd68312;
    data[3709] = -'sd69390;
    data[3710] =  'sd67501;
    data[3711] =  'sd49115;
    data[3712] =  'sd80988;
    data[3713] =  'sd58608;
    data[3714] = -'sd9369;
    data[3715] = -'sd70384;
    data[3716] =  'sd42651;
    data[3717] = -'sd80612;
    data[3718] = -'sd49208;
    data[3719] =  'sd80528;
    data[3720] =  'sd47108;
    data[3721] =  'sd30813;
    data[3722] = -'sd48880;
    data[3723] = -'sd75113;
    data[3724] = -'sd75574;
    data[3725] =  'sd76742;
    data[3726] = -'sd47542;
    data[3727] = -'sd41663;
    data[3728] = -'sd58529;
    data[3729] =  'sd11344;
    data[3730] = -'sd44082;
    data[3731] =  'sd44837;
    data[3732] = -'sd25962;
    data[3733] =  'sd6314;
    data[3734] = -'sd5991;
    data[3735] =  'sd14066;
    data[3736] =  'sd23968;
    data[3737] = -'sd56164;
    data[3738] =  'sd70469;
    data[3739] = -'sd40526;
    data[3740] = -'sd30104;
    data[3741] =  'sd66605;
    data[3742] =  'sd26715;
    data[3743] =  'sd12511;
    data[3744] = -'sd14907;
    data[3745] = -'sd44993;
    data[3746] =  'sd22062;
    data[3747] =  'sd60027;
    data[3748] =  'sd26106;
    data[3749] = -'sd2714;
    data[3750] = -'sd67850;
    data[3751] = -'sd57840;
    data[3752] =  'sd28569;
    data[3753] =  'sd58861;
    data[3754] = -'sd3044;
    data[3755] = -'sd76100;
    data[3756] =  'sd63592;
    data[3757] = -'sd48610;
    data[3758] = -'sd68363;
    data[3759] = -'sd70665;
    data[3760] =  'sd35626;
    data[3761] =  'sd71445;
    data[3762] = -'sd16126;
    data[3763] = -'sd75468;
    data[3764] =  'sd79392;
    data[3765] =  'sd18708;
    data[3766] = -'sd23823;
    data[3767] =  'sd59789;
    data[3768] =  'sd20156;
    data[3769] =  'sd12377;
    data[3770] = -'sd18257;
    data[3771] =  'sd35098;
    data[3772] =  'sd58245;
    data[3773] = -'sd18444;
    data[3774] =  'sd30423;
    data[3775] = -'sd58630;
    data[3776] =  'sd8819;
    data[3777] =  'sd56634;
    data[3778] = -'sd58719;
    data[3779] =  'sd6594;
    data[3780] =  'sd1009;
    data[3781] =  'sd25225;
    data[3782] = -'sd24739;
    data[3783] =  'sd36889;
    data[3784] = -'sd60821;
    data[3785] = -'sd45956;
    data[3786] = -'sd2013;
    data[3787] = -'sd50325;
    data[3788] =  'sd52603;
    data[3789] =  'sd4347;
    data[3790] = -'sd55166;
    data[3791] = -'sd68422;
    data[3792] = -'sd72140;
    data[3793] = -'sd1249;
    data[3794] = -'sd31225;
    data[3795] =  'sd38580;
    data[3796] = -'sd18546;
    data[3797] =  'sd27873;
    data[3798] =  'sd41461;
    data[3799] =  'sd53479;
    data[3800] =  'sd26247;
    data[3801] =  'sd811;
    data[3802] =  'sd20275;
    data[3803] =  'sd15352;
    data[3804] =  'sd56118;
    data[3805] = -'sd71619;
    data[3806] =  'sd11776;
    data[3807] = -'sd33282;
    data[3808] = -'sd12845;
    data[3809] =  'sd6557;
    data[3810] =  'sd84;
    data[3811] =  'sd2100;
    data[3812] =  'sd52500;
    data[3813] =  'sd1772;
    data[3814] =  'sd44300;
    data[3815] = -'sd39387;
    data[3816] = -'sd1629;
    data[3817] = -'sd40725;
    data[3818] = -'sd35079;
    data[3819] = -'sd57770;
    data[3820] =  'sd30319;
    data[3821] = -'sd61230;
    data[3822] = -'sd56181;
    data[3823] =  'sd70044;
    data[3824] = -'sd51151;
    data[3825] =  'sd31953;
    data[3826] = -'sd20380;
    data[3827] = -'sd17977;
    data[3828] =  'sd42098;
    data[3829] =  'sd69404;
    data[3830] = -'sd67151;
    data[3831] = -'sd40365;
    data[3832] = -'sd26079;
    data[3833] =  'sd3389;
    data[3834] = -'sd79116;
    data[3835] = -'sd11808;
    data[3836] =  'sd32482;
    data[3837] = -'sd7155;
    data[3838] = -'sd15034;
    data[3839] = -'sd48168;
    data[3840] = -'sd57313;
    data[3841] =  'sd41744;
    data[3842] =  'sd60554;
    data[3843] =  'sd39281;
    data[3844] = -'sd1021;
    data[3845] = -'sd25525;
    data[3846] =  'sd17239;
    data[3847] = -'sd60548;
    data[3848] = -'sd39131;
    data[3849] =  'sd4771;
    data[3850] = -'sd44566;
    data[3851] =  'sd32737;
    data[3852] = -'sd780;
    data[3853] = -'sd19500;
    data[3854] =  'sd4023;
    data[3855] = -'sd63266;
    data[3856] =  'sd56760;
    data[3857] = -'sd55569;
    data[3858] = -'sd78497;
    data[3859] =  'sd3667;
    data[3860] = -'sd72166;
    data[3861] = -'sd1899;
    data[3862] = -'sd47475;
    data[3863] = -'sd39988;
    data[3864] = -'sd16654;
    data[3865] =  'sd75173;
    data[3866] =  'sd77074;
    data[3867] = -'sd39242;
    data[3868] =  'sd1996;
    data[3869] =  'sd49900;
    data[3870] = -'sd63228;
    data[3871] =  'sd57710;
    data[3872] = -'sd31819;
    data[3873] =  'sd23730;
    data[3874] = -'sd62114;
    data[3875] = -'sd78281;
    data[3876] =  'sd9067;
    data[3877] =  'sd62834;
    data[3878] = -'sd67560;
    data[3879] = -'sd50590;
    data[3880] =  'sd45978;
    data[3881] =  'sd2563;
    data[3882] =  'sd64075;
    data[3883] = -'sd36535;
    data[3884] =  'sd69671;
    data[3885] = -'sd60476;
    data[3886] = -'sd37331;
    data[3887] =  'sd49771;
    data[3888] = -'sd66453;
    data[3889] = -'sd22915;
    data[3890] = -'sd81352;
    data[3891] = -'sd67708;
    data[3892] = -'sd54290;
    data[3893] = -'sd46522;
    data[3894] = -'sd16163;
    data[3895] = -'sd76393;
    data[3896] =  'sd56267;
    data[3897] = -'sd67894;
    data[3898] = -'sd58940;
    data[3899] =  'sd1069;
    data[3900] =  'sd26725;
    data[3901] =  'sd12761;
    data[3902] = -'sd8657;
    data[3903] = -'sd52584;
    data[3904] = -'sd3872;
    data[3905] =  'sd67041;
    data[3906] =  'sd37615;
    data[3907] = -'sd42671;
    data[3908] =  'sd80112;
    data[3909] =  'sd36708;
    data[3910] = -'sd65346;
    data[3911] =  'sd4760;
    data[3912] = -'sd44841;
    data[3913] =  'sd25862;
    data[3914] = -'sd8814;
    data[3915] = -'sd56509;
    data[3916] =  'sd61844;
    data[3917] =  'sd71531;
    data[3918] = -'sd13976;
    data[3919] = -'sd21718;
    data[3920] = -'sd51427;
    data[3921] =  'sd25053;
    data[3922] = -'sd29039;
    data[3923] = -'sd70611;
    data[3924] =  'sd36976;
    data[3925] = -'sd58646;
    data[3926] =  'sd8419;
    data[3927] =  'sd46634;
    data[3928] =  'sd18963;
    data[3929] = -'sd17448;
    data[3930] =  'sd55323;
    data[3931] =  'sd72347;
    data[3932] =  'sd6424;
    data[3933] = -'sd3241;
    data[3934] = -'sd81025;
    data[3935] = -'sd59533;
    data[3936] = -'sd13756;
    data[3937] = -'sd16218;
    data[3938] = -'sd77768;
    data[3939] =  'sd21892;
    data[3940] =  'sd55777;
    data[3941] = -'sd80144;
    data[3942] = -'sd37508;
    data[3943] =  'sd45346;
    data[3944] = -'sd13237;
    data[3945] = -'sd3243;
    data[3946] = -'sd81075;
    data[3947] = -'sd60783;
    data[3948] = -'sd45006;
    data[3949] =  'sd21737;
    data[3950] =  'sd51902;
    data[3951] = -'sd13178;
    data[3952] = -'sd1768;
    data[3953] = -'sd44200;
    data[3954] =  'sd41887;
    data[3955] =  'sd64129;
    data[3956] = -'sd35185;
    data[3957] = -'sd60420;
    data[3958] = -'sd35931;
    data[3959] = -'sd79070;
    data[3960] = -'sd10658;
    data[3961] =  'sd61232;
    data[3962] =  'sd56231;
    data[3963] = -'sd68794;
    data[3964] = -'sd81440;
    data[3965] = -'sd69908;
    data[3966] =  'sd54551;
    data[3967] =  'sd53047;
    data[3968] =  'sd15447;
    data[3969] =  'sd58493;
    data[3970] = -'sd12244;
    data[3971] =  'sd21582;
    data[3972] =  'sd48027;
    data[3973] =  'sd53788;
    data[3974] =  'sd33972;
    data[3975] =  'sd30095;
    data[3976] = -'sd66830;
    data[3977] = -'sd32340;
    data[3978] =  'sd10705;
    data[3979] = -'sd60057;
    data[3980] = -'sd26856;
    data[3981] = -'sd16036;
    data[3982] = -'sd73218;
    data[3983] = -'sd28199;
    data[3984] = -'sd49611;
    data[3985] =  'sd70453;
    data[3986] = -'sd40926;
    data[3987] = -'sd40104;
    data[3988] = -'sd19554;
    data[3989] =  'sd2673;
    data[3990] =  'sd66825;
    data[3991] =  'sd32215;
    data[3992] = -'sd13830;
    data[3993] = -'sd18068;
    data[3994] =  'sd39823;
    data[3995] =  'sd12529;
    data[3996] = -'sd14457;
    data[3997] = -'sd33743;
    data[3998] = -'sd24370;
    data[3999] =  'sd46114;
    data[4000] =  'sd5963;
    data[4001] = -'sd14766;
    data[4002] = -'sd41468;
    data[4003] = -'sd53654;
    data[4004] = -'sd30622;
    data[4005] =  'sd53655;
    data[4006] =  'sd30647;
    data[4007] = -'sd53030;
    data[4008] = -'sd15022;
    data[4009] = -'sd47868;
    data[4010] = -'sd49813;
    data[4011] =  'sd65403;
    data[4012] = -'sd3335;
    data[4013] =  'sd80466;
    data[4014] =  'sd45558;
    data[4015] = -'sd7937;
    data[4016] = -'sd34584;
    data[4017] = -'sd45395;
    data[4018] =  'sd12012;
    data[4019] = -'sd27382;
    data[4020] = -'sd29186;
    data[4021] = -'sd74286;
    data[4022] = -'sd54899;
    data[4023] = -'sd61747;
    data[4024] = -'sd69106;
    data[4025] =  'sd74601;
    data[4026] =  'sd62774;
    data[4027] = -'sd69060;
    data[4028] =  'sd75751;
    data[4029] = -'sd72317;
    data[4030] = -'sd5674;
    data[4031] =  'sd21991;
    data[4032] =  'sd58252;
    data[4033] = -'sd18269;
    data[4034] =  'sd34798;
    data[4035] =  'sd50745;
    data[4036] = -'sd42103;
    data[4037] = -'sd69529;
    data[4038] =  'sd64026;
    data[4039] = -'sd37760;
    data[4040] =  'sd39046;
    data[4041] = -'sd6896;
    data[4042] = -'sd8559;
    data[4043] = -'sd50134;
    data[4044] =  'sd57378;
    data[4045] = -'sd40119;
    data[4046] = -'sd19929;
    data[4047] = -'sd6702;
    data[4048] = -'sd3709;
    data[4049] =  'sd71116;
    data[4050] = -'sd24351;
    data[4051] =  'sd46589;
    data[4052] =  'sd17838;
    data[4053] = -'sd45573;
    data[4054] =  'sd7562;
    data[4055] =  'sd25209;
    data[4056] = -'sd25139;
    data[4057] =  'sd26889;
    data[4058] =  'sd16861;
    data[4059] = -'sd69998;
    data[4060] =  'sd52301;
    data[4061] = -'sd3203;
    data[4062] = -'sd80075;
    data[4063] = -'sd35783;
    data[4064] = -'sd75370;
    data[4065] =  'sd81842;
    data[4066] =  'sd79958;
    data[4067] =  'sd32858;
    data[4068] =  'sd2245;
    data[4069] =  'sd56125;
    data[4070] = -'sd71444;
    data[4071] =  'sd16151;
    data[4072] =  'sd76093;
    data[4073] = -'sd63767;
    data[4074] =  'sd44235;
    data[4075] = -'sd41012;
    data[4076] = -'sd42254;
    data[4077] = -'sd73304;
    data[4078] = -'sd30349;
    data[4079] =  'sd60480;
    data[4080] =  'sd37431;
    data[4081] = -'sd47271;
    data[4082] = -'sd34888;
    data[4083] = -'sd52995;
    data[4084] = -'sd14147;
    data[4085] = -'sd25993;
    data[4086] =  'sd5539;
    data[4087] = -'sd25366;
    data[4088] =  'sd21214;
    data[4089] =  'sd38827;
    data[4090] = -'sd12371;
    data[4091] =  'sd18407;
    data[4092] = -'sd31348;
    data[4093] =  'sd35505;
    data[4094] =  'sd68420;
    data[4095] =  'sd72090;
  end

endmodule

