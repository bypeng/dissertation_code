module f_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [12:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd1195; // 0
        'h001: dout <= -'sd1779; // 1
        'h002: dout <= -'sd206; // 2
        'h003: dout <= -'sd1330; // 3
        'h004: dout <=  'sd1763; // 4
        'h005: dout <=  'sd1387; // 5
        'h006: dout <=  'sd1573; // 6
        'h007: dout <=  'sd814; // 7
        'h008: dout <= -'sd576; // 8
        'h009: dout <= -'sd1527; // 9
        'h00a: dout <=  'sd1701; // 10
        'h00b: dout <= -'sd2063; // 11
        'h00c: dout <=  'sd898; // 12
        'h00d: dout <=  'sd1250; // 13
        'h00e: dout <= -'sd2278; // 14
        'h00f: dout <=  'sd1353; // 15
        'h010: dout <= -'sd114; // 16
        'h011: dout <= -'sd421; // 17
        'h012: dout <= -'sd1458; // 18
        'h013: dout <=  'sd305; // 19
        'h014: dout <= -'sd2045; // 20
        'h015: dout <= -'sd2113; // 21
        'h016: dout <= -'sd2087; // 22
        'h017: dout <=  'sd2140; // 23
        'h018: dout <= -'sd2220; // 24
        'h019: dout <=  'sd827; // 25
        'h01a: dout <= -'sd521; // 26
        'h01b: dout <=  'sd1162; // 27
        'h01c: dout <= -'sd2058; // 28
        'h01d: dout <=  'sd2027; // 29
        'h01e: dout <= -'sd479; // 30
        'h01f: dout <=  'sd1292; // 31
        'h020: dout <=  'sd1766; // 32
        'h021: dout <=  'sd2234; // 33
        'h022: dout <= -'sd386; // 34
        'h023: dout <=  'sd536; // 35
        'h024: dout <= -'sd404; // 36
        'h025: dout <= -'sd503; // 37
        'h026: dout <=  'sd1470; // 38
        'h027: dout <=  'sd78; // 39
        'h028: dout <= -'sd2119; // 40
        'h029: dout <=  'sd1114; // 41
        'h02a: dout <=  'sd2263; // 42
        'h02b: dout <= -'sd1476; // 43
        'h02c: dout <= -'sd773; // 44
        'h02d: dout <=  'sd133; // 45
        'h02e: dout <= -'sd1305; // 46
        'h02f: dout <=  'sd430; // 47
        'h030: dout <=  'sd1807; // 48
        'h031: dout <=  'sd1162; // 49
        'h032: dout <=  'sd1864; // 50
        'h033: dout <= -'sd740; // 51
        'h034: dout <=  'sd190; // 52
        'h035: dout <=  'sd32; // 53
        'h036: dout <=  'sd1795; // 54
        'h037: dout <=  'sd1844; // 55
        'h038: dout <=  'sd927; // 56
        'h039: dout <= -'sd2013; // 57
        'h03a: dout <=  'sd1639; // 58
        'h03b: dout <= -'sd307; // 59
        'h03c: dout <=  'sd1016; // 60
        'h03d: dout <=  'sd1099; // 61
        'h03e: dout <= -'sd878; // 62
        'h03f: dout <=  'sd712; // 63
        'h040: dout <=  'sd2200; // 64
        'h041: dout <=  'sd774; // 65
        'h042: dout <= -'sd1587; // 66
        'h043: dout <=  'sd1300; // 67
        'h044: dout <=  'sd1870; // 68
        'h045: dout <= -'sd1411; // 69
        'h046: dout <= -'sd954; // 70
        'h047: dout <=  'sd1972; // 71
        'h048: dout <=  'sd926; // 72
        'h049: dout <=  'sd740; // 73
        'h04a: dout <=  'sd1716; // 74
        'h04b: dout <= -'sd2053; // 75
        'h04c: dout <=  'sd1549; // 76
        'h04d: dout <= -'sd1939; // 77
        'h04e: dout <=  'sd232; // 78
        'h04f: dout <=  'sd929; // 79
        'h050: dout <= -'sd900; // 80
        'h051: dout <= -'sd914; // 81
        'h052: dout <=  'sd1819; // 82
        'h053: dout <= -'sd436; // 83
        'h054: dout <= -'sd2195; // 84
        'h055: dout <= -'sd661; // 85
        'h056: dout <=  'sd2125; // 86
        'h057: dout <=  'sd2196; // 87
        'h058: dout <= -'sd394; // 88
        'h059: dout <=  'sd1018; // 89
        'h05a: dout <=  'sd1913; // 90
        'h05b: dout <=  'sd521; // 91
        'h05c: dout <=  'sd599; // 92
        'h05d: dout <=  'sd1466; // 93
        'h05e: dout <= -'sd90; // 94
        'h05f: dout <=  'sd2194; // 95
        'h060: dout <= -'sd2249; // 96
        'h061: dout <=  'sd848; // 97
        'h062: dout <=  'sd1903; // 98
        'h063: dout <= -'sd1237; // 99
        'h064: dout <=  'sd1954; // 100
        'h065: dout <= -'sd612; // 101
        'h066: dout <=  'sd1195; // 102
        'h067: dout <= -'sd1836; // 103
        'h068: dout <=  'sd1646; // 104
        'h069: dout <=  'sd692; // 105
        'h06a: dout <=  'sd2246; // 106
        'h06b: dout <= -'sd658; // 107
        'h06c: dout <=  'sd1839; // 108
        'h06d: dout <=  'sd1091; // 109
        'h06e: dout <=  'sd1677; // 110
        'h06f: dout <=  'sd627; // 111
        'h070: dout <=  'sd1099; // 112
        'h071: dout <=  'sd540; // 113
        'h072: dout <= -'sd2283; // 114
        'h073: dout <=  'sd2116; // 115
        'h074: dout <=  'sd2129; // 116
        'h075: dout <=  'sd417; // 117
        'h076: dout <=  'sd1458; // 118
        'h077: dout <= -'sd2066; // 119
        'h078: dout <= -'sd415; // 120
        'h079: dout <= -'sd844; // 121
        'h07a: dout <=  'sd2216; // 122
        'h07b: dout <= -'sd815; // 123
        'h07c: dout <= -'sd1545; // 124
        'h07d: dout <=  'sd2219; // 125
        'h07e: dout <= -'sd204; // 126
        'h07f: dout <= -'sd2030; // 127
        'h080: dout <= -'sd1718; // 128
        'h081: dout <= -'sd1614; // 129
        'h082: dout <= -'sd2159; // 130
        'h083: dout <=  'sd1415; // 131
        'h084: dout <= -'sd2176; // 132
        'h085: dout <=  'sd8; // 133
        'h086: dout <= -'sd251; // 134
        'h087: dout <= -'sd95; // 135
        'h088: dout <= -'sd1399; // 136
        'h089: dout <= -'sd783; // 137
        'h08a: dout <=  'sd526; // 138
        'h08b: dout <=  'sd83; // 139
        'h08c: dout <= -'sd1726; // 140
        'h08d: dout <= -'sd924; // 141
        'h08e: dout <= -'sd988; // 142
        'h08f: dout <= -'sd205; // 143
        'h090: dout <=  'sd2025; // 144
        'h091: dout <= -'sd918; // 145
        'h092: dout <= -'sd60; // 146
        'h093: dout <=  'sd117; // 147
        'h094: dout <=  'sd1429; // 148
        'h095: dout <=  'sd342; // 149
        'h096: dout <=  'sd1772; // 150
        'h097: dout <=  'sd1586; // 151
        'h098: dout <= -'sd1360; // 152
        'h099: dout <= -'sd2102; // 153
        'h09a: dout <=  'sd260; // 154
        'h09b: dout <=  'sd871; // 155
        'h09c: dout <=  'sd517; // 156
        'h09d: dout <=  'sd1153; // 157
        'h09e: dout <= -'sd755; // 158
        'h09f: dout <= -'sd179; // 159
        'h0a0: dout <= -'sd1405; // 160
        'h0a1: dout <= -'sd219; // 161
        'h0a2: dout <=  'sd1883; // 162
        'h0a3: dout <= -'sd583; // 163
        'h0a4: dout <=  'sd1241; // 164
        'h0a5: dout <= -'sd2125; // 165
        'h0a6: dout <= -'sd449; // 166
        'h0a7: dout <= -'sd2149; // 167
        'h0a8: dout <=  'sd959; // 168
        'h0a9: dout <= -'sd1096; // 169
        'h0aa: dout <= -'sd2006; // 170
        'h0ab: dout <= -'sd983; // 171
        'h0ac: dout <=  'sd1355; // 172
        'h0ad: dout <=  'sd1852; // 173
        'h0ae: dout <=  'sd1200; // 174
        'h0af: dout <=  'sd2167; // 175
        'h0b0: dout <= -'sd488; // 176
        'h0b1: dout <=  'sd1936; // 177
        'h0b2: dout <=  'sd1398; // 178
        'h0b3: dout <= -'sd467; // 179
        'h0b4: dout <=  'sd1996; // 180
        'h0b5: dout <= -'sd2044; // 181
        'h0b6: dout <=  'sd940; // 182
        'h0b7: dout <=  'sd336; // 183
        'h0b8: dout <=  'sd1197; // 184
        'h0b9: dout <= -'sd1814; // 185
        'h0ba: dout <=  'sd151; // 186
        'h0bb: dout <= -'sd1266; // 187
        'h0bc: dout <= -'sd558; // 188
        'h0bd: dout <= -'sd1907; // 189
        'h0be: dout <=  'sd214; // 190
        'h0bf: dout <= -'sd1716; // 191
        'h0c0: dout <= -'sd1669; // 192
        'h0c1: dout <=  'sd247; // 193
        'h0c2: dout <=  'sd145; // 194
        'h0c3: dout <= -'sd999; // 195
        'h0c4: dout <=  'sd1114; // 196
        'h0c5: dout <= -'sd228; // 197
        'h0c6: dout <= -'sd1227; // 198
        'h0c7: dout <= -'sd2226; // 199
        'h0c8: dout <= -'sd1985; // 200
        'h0c9: dout <= -'sd513; // 201
        'h0ca: dout <=  'sd1480; // 202
        'h0cb: dout <= -'sd890; // 203
        'h0cc: dout <=  'sd1873; // 204
        'h0cd: dout <= -'sd1989; // 205
        'h0ce: dout <=  'sd801; // 206
        'h0cf: dout <= -'sd654; // 207
        'h0d0: dout <=  'sd547; // 208
        'h0d1: dout <= -'sd1484; // 209
        'h0d2: dout <= -'sd610; // 210
        'h0d3: dout <=  'sd1251; // 211
        'h0d4: dout <= -'sd705; // 212
        'h0d5: dout <=  'sd1738; // 213
        'h0d6: dout <= -'sd1440; // 214
        'h0d7: dout <=  'sd900; // 215
        'h0d8: dout <=  'sd130; // 216
        'h0d9: dout <=  'sd1834; // 217
        'h0da: dout <=  'sd1799; // 218
        'h0db: dout <= -'sd2155; // 219
        'h0dc: dout <=  'sd370; // 220
        'h0dd: dout <=  'sd1000; // 221
        'h0de: dout <=  'sd9; // 222
        'h0df: dout <= -'sd2147; // 223
        'h0e0: dout <= -'sd1010; // 224
        'h0e1: dout <= -'sd650; // 225
        'h0e2: dout <=  'sd389; // 226
        'h0e3: dout <= -'sd1188; // 227
        'h0e4: dout <=  'sd482; // 228
        'h0e5: dout <=  'sd1221; // 229
        'h0e6: dout <= -'sd550; // 230
        'h0e7: dout <= -'sd112; // 231
        'h0e8: dout <= -'sd1506; // 232
        'h0e9: dout <=  'sd811; // 233
        'h0ea: dout <=  'sd2191; // 234
        'h0eb: dout <=  'sd521; // 235
        'h0ec: dout <=  'sd2082; // 236
        'h0ed: dout <=  'sd1674; // 237
        'h0ee: dout <=  'sd2067; // 238
        'h0ef: dout <= -'sd373; // 239
        'h0f0: dout <= -'sd1760; // 240
        'h0f1: dout <= -'sd1965; // 241
        'h0f2: dout <= -'sd1602; // 242
        'h0f3: dout <= -'sd1206; // 243
        'h0f4: dout <= -'sd905; // 244
        'h0f5: dout <= -'sd931; // 245
        'h0f6: dout <=  'sd2114; // 246
        'h0f7: dout <= -'sd551; // 247
        'h0f8: dout <= -'sd100; // 248
        'h0f9: dout <=  'sd426; // 249
        'h0fa: dout <=  'sd1849; // 250
        'h0fb: dout <= -'sd204; // 251
        'h0fc: dout <=  'sd720; // 252
        'h0fd: dout <=  'sd480; // 253
        'h0fe: dout <=  'sd492; // 254
        'h0ff: dout <= -'sd1362; // 255
        'h100: dout <=  'sd90; // 256
        'h101: dout <= -'sd369; // 257
        'h102: dout <=  'sd1709; // 258
        'h103: dout <= -'sd1187; // 259
        'h104: dout <=  'sd2220; // 260
        'h105: dout <= -'sd1441; // 261
        'h106: dout <=  'sd332; // 262
        'h107: dout <= -'sd1975; // 263
        'h108: dout <=  'sd1035; // 264
        'h109: dout <= -'sd1696; // 265
        'h10a: dout <=  'sd819; // 266
        'h10b: dout <= -'sd1089; // 267
        'h10c: dout <= -'sd1271; // 268
        'h10d: dout <=  'sd497; // 269
        'h10e: dout <= -'sd1356; // 270
        'h10f: dout <=  'sd801; // 271
        'h110: dout <= -'sd1668; // 272
        'h111: dout <=  'sd2212; // 273
        'h112: dout <= -'sd463; // 274
        'h113: dout <= -'sd1626; // 275
        'h114: dout <= -'sd110; // 276
        'h115: dout <=  'sd694; // 277
        'h116: dout <=  'sd126; // 278
        'h117: dout <=  'sd2081; // 279
        'h118: dout <= -'sd1359; // 280
        'h119: dout <=  'sd1455; // 281
        'h11a: dout <= -'sd25; // 282
        'h11b: dout <= -'sd1413; // 283
        'h11c: dout <= -'sd1921; // 284
        'h11d: dout <=  'sd127; // 285
        'h11e: dout <= -'sd2194; // 286
        'h11f: dout <= -'sd2176; // 287
        'h120: dout <= -'sd1544; // 288
        'h121: dout <=  'sd1092; // 289
        'h122: dout <= -'sd1353; // 290
        'h123: dout <= -'sd1968; // 291
        'h124: dout <= -'sd756; // 292
        'h125: dout <= -'sd332; // 293
        'h126: dout <=  'sd1153; // 294
        'h127: dout <= -'sd968; // 295
        'h128: dout <= -'sd1349; // 296
        'h129: dout <=  'sd1398; // 297
        'h12a: dout <= -'sd924; // 298
        'h12b: dout <= -'sd318; // 299
        'h12c: dout <= -'sd993; // 300
        'h12d: dout <= -'sd1453; // 301
        'h12e: dout <=  'sd1269; // 302
        'h12f: dout <=  'sd803; // 303
        'h130: dout <=  'sd2152; // 304
        'h131: dout <=  'sd113; // 305
        'h132: dout <=  'sd2212; // 306
        'h133: dout <= -'sd220; // 307
        'h134: dout <=  'sd1612; // 308
        'h135: dout <=  'sd281; // 309
        'h136: dout <= -'sd1475; // 310
        'h137: dout <= -'sd595; // 311
        'h138: dout <=  'sd305; // 312
        'h139: dout <= -'sd1971; // 313
        'h13a: dout <= -'sd2072; // 314
        'h13b: dout <= -'sd2209; // 315
        'h13c: dout <=  'sd126; // 316
        'h13d: dout <=  'sd328; // 317
        'h13e: dout <=  'sd1390; // 318
        'h13f: dout <=  'sd910; // 319
        'h140: dout <=  'sd271; // 320
        'h141: dout <=  'sd969; // 321
        'h142: dout <= -'sd1780; // 322
        'h143: dout <= -'sd1770; // 323
        'h144: dout <=  'sd304; // 324
        'h145: dout <=  'sd1439; // 325
        'h146: dout <= -'sd1383; // 326
        'h147: dout <= -'sd247; // 327
        'h148: dout <= -'sd533; // 328
        'h149: dout <=  'sd2152; // 329
        'h14a: dout <=  'sd1546; // 330
        'h14b: dout <=  'sd619; // 331
        'h14c: dout <= -'sd173; // 332
        'h14d: dout <= -'sd795; // 333
        'h14e: dout <=  'sd2141; // 334
        'h14f: dout <= -'sd593; // 335
        'h150: dout <=  'sd222; // 336
        'h151: dout <= -'sd664; // 337
        'h152: dout <= -'sd277; // 338
        'h153: dout <=  'sd657; // 339
        'h154: dout <= -'sd1629; // 340
        'h155: dout <=  'sd5; // 341
        'h156: dout <= -'sd1563; // 342
        'h157: dout <=  'sd1374; // 343
        'h158: dout <= -'sd1554; // 344
        'h159: dout <=  'sd481; // 345
        'h15a: dout <= -'sd432; // 346
        'h15b: dout <=  'sd903; // 347
        'h15c: dout <=  'sd218; // 348
        'h15d: dout <= -'sd1959; // 349
        'h15e: dout <=  'sd385; // 350
        'h15f: dout <= -'sd765; // 351
        'h160: dout <=  'sd299; // 352
        'h161: dout <=  'sd185; // 353
        'h162: dout <= -'sd282; // 354
        'h163: dout <=  'sd443; // 355
        'h164: dout <= -'sd1469; // 356
        'h165: dout <=  'sd2163; // 357
        'h166: dout <= -'sd1541; // 358
        'h167: dout <= -'sd288; // 359
        'h168: dout <= -'sd492; // 360
        'h169: dout <= -'sd2129; // 361
        'h16a: dout <= -'sd299; // 362
        'h16b: dout <=  'sd996; // 363
        'h16c: dout <= -'sd1703; // 364
        'h16d: dout <= -'sd100; // 365
        'h16e: dout <=  'sd2220; // 366
        'h16f: dout <= -'sd1715; // 367
        'h170: dout <= -'sd1680; // 368
        'h171: dout <= -'sd2119; // 369
        'h172: dout <= -'sd2214; // 370
        'h173: dout <=  'sd87; // 371
        'h174: dout <=  'sd647; // 372
        'h175: dout <=  'sd1745; // 373
        'h176: dout <=  'sd1545; // 374
        'h177: dout <= -'sd1032; // 375
        'h178: dout <= -'sd1469; // 376
        'h179: dout <=  'sd1812; // 377
        'h17a: dout <=  'sd392; // 378
        'h17b: dout <= -'sd1664; // 379
        'h17c: dout <=  'sd1876; // 380
        'h17d: dout <= -'sd876; // 381
        'h17e: dout <= -'sd824; // 382
        'h17f: dout <= -'sd1070; // 383
        'h180: dout <= -'sd1136; // 384
        'h181: dout <=  'sd324; // 385
        'h182: dout <=  'sd208; // 386
        'h183: dout <= -'sd1420; // 387
        'h184: dout <=  'sd1918; // 388
        'h185: dout <=  'sd109; // 389
        'h186: dout <= -'sd1261; // 390
        'h187: dout <= -'sd602; // 391
        'h188: dout <= -'sd1135; // 392
        'h189: dout <=  'sd2173; // 393
        'h18a: dout <= -'sd2035; // 394
        'h18b: dout <=  'sd294; // 395
        'h18c: dout <=  'sd2234; // 396
        'h18d: dout <= -'sd613; // 397
        'h18e: dout <= -'sd836; // 398
        'h18f: dout <=  'sd153; // 399
        'h190: dout <=  'sd1249; // 400
        'h191: dout <=  'sd2108; // 401
        'h192: dout <= -'sd1002; // 402
        'h193: dout <= -'sd1898; // 403
        'h194: dout <= -'sd270; // 404
        'h195: dout <= -'sd226; // 405
        'h196: dout <= -'sd1768; // 406
        'h197: dout <=  'sd1364; // 407
        'h198: dout <=  'sd1228; // 408
        'h199: dout <=  'sd2204; // 409
        'h19a: dout <= -'sd246; // 410
        'h19b: dout <=  'sd2139; // 411
        'h19c: dout <=  'sd1304; // 412
        'h19d: dout <=  'sd2112; // 413
        'h19e: dout <=  'sd1418; // 414
        'h19f: dout <= -'sd2206; // 415
        'h1a0: dout <=  'sd946; // 416
        'h1a1: dout <=  'sd479; // 417
        'h1a2: dout <= -'sd890; // 418
        'h1a3: dout <= -'sd182; // 419
        'h1a4: dout <=  'sd1684; // 420
        'h1a5: dout <= -'sd2096; // 421
        'h1a6: dout <=  'sd1118; // 422
        'h1a7: dout <= -'sd2141; // 423
        'h1a8: dout <= -'sd1785; // 424
        'h1a9: dout <=  'sd612; // 425
        'h1aa: dout <= -'sd1163; // 426
        'h1ab: dout <= -'sd1270; // 427
        'h1ac: dout <= -'sd1161; // 428
        'h1ad: dout <= -'sd173; // 429
        'h1ae: dout <= -'sd27; // 430
        'h1af: dout <=  'sd963; // 431
        'h1b0: dout <=  'sd990; // 432
        'h1b1: dout <= -'sd885; // 433
        'h1b2: dout <= -'sd1564; // 434
        'h1b3: dout <= -'sd382; // 435
        'h1b4: dout <=  'sd1686; // 436
        'h1b5: dout <= -'sd2234; // 437
        'h1b6: dout <= -'sd841; // 438
        'h1b7: dout <=  'sd2036; // 439
        'h1b8: dout <=  'sd303; // 440
        'h1b9: dout <=  'sd1808; // 441
        'h1ba: dout <=  'sd1295; // 442
        'h1bb: dout <= -'sd446; // 443
        'h1bc: dout <= -'sd343; // 444
        'h1bd: dout <=  'sd268; // 445
        'h1be: dout <=  'sd1760; // 446
        'h1bf: dout <=  'sd1627; // 447
        'h1c0: dout <= -'sd452; // 448
        'h1c1: dout <=  'sd1082; // 449
        'h1c2: dout <=  'sd465; // 450
        'h1c3: dout <=  'sd2295; // 451
        'h1c4: dout <= -'sd41; // 452
        'h1c5: dout <= -'sd498; // 453
        'h1c6: dout <= -'sd1901; // 454
        'h1c7: dout <= -'sd1709; // 455
        'h1c8: dout <=  'sd1896; // 456
        'h1c9: dout <=  'sd725; // 457
        'h1ca: dout <= -'sd989; // 458
        'h1cb: dout <=  'sd1896; // 459
        'h1cc: dout <= -'sd626; // 460
        'h1cd: dout <=  'sd259; // 461
        'h1ce: dout <=  'sd152; // 462
        'h1cf: dout <=  'sd159; // 463
        'h1d0: dout <=  'sd2229; // 464
        'h1d1: dout <=  'sd749; // 465
        'h1d2: dout <= -'sd942; // 466
        'h1d3: dout <=  'sd1512; // 467
        'h1d4: dout <= -'sd1599; // 468
        'h1d5: dout <= -'sd1286; // 469
        'h1d6: dout <=  'sd1915; // 470
        'h1d7: dout <=  'sd795; // 471
        'h1d8: dout <= -'sd851; // 472
        'h1d9: dout <= -'sd1019; // 473
        'h1da: dout <= -'sd243; // 474
        'h1db: dout <=  'sd1200; // 475
        'h1dc: dout <= -'sd513; // 476
        'h1dd: dout <= -'sd1868; // 477
        'h1de: dout <=  'sd1760; // 478
        'h1df: dout <=  'sd929; // 479
        'h1e0: dout <=  'sd555; // 480
        'h1e1: dout <=  'sd850; // 481
        'h1e2: dout <=  'sd1924; // 482
        'h1e3: dout <= -'sd945; // 483
        'h1e4: dout <=  'sd2163; // 484
        'h1e5: dout <= -'sd1962; // 485
        'h1e6: dout <=  'sd1999; // 486
        'h1e7: dout <= -'sd1555; // 487
        'h1e8: dout <= -'sd205; // 488
        'h1e9: dout <= -'sd1468; // 489
        'h1ea: dout <= -'sd104; // 490
        'h1eb: dout <= -'sd1610; // 491
        'h1ec: dout <= -'sd1156; // 492
        'h1ed: dout <= -'sd1624; // 493
        'h1ee: dout <=  'sd1350; // 494
        'h1ef: dout <= -'sd321; // 495
        'h1f0: dout <=  'sd837; // 496
        'h1f1: dout <=  'sd1251; // 497
        'h1f2: dout <=  'sd959; // 498
        'h1f3: dout <= -'sd946; // 499
        'h1f4: dout <=  'sd371; // 500
        'h1f5: dout <=  'sd1294; // 501
        'h1f6: dout <= -'sd1261; // 502
        'h1f7: dout <=  'sd1702; // 503
        'h1f8: dout <= -'sd559; // 504
        'h1f9: dout <= -'sd1319; // 505
        'h1fa: dout <=  'sd1237; // 506
        'h1fb: dout <=  'sd2079; // 507
        'h1fc: dout <=  'sd1049; // 508
        'h1fd: dout <= -'sd1328; // 509
        'h1fe: dout <=  'sd125; // 510
        'h1ff: dout <= -'sd21; // 511
        'h200: dout <= -'sd262; // 512
        'h201: dout <=  'sd808; // 513
        'h202: dout <=  'sd2287; // 514
        'h203: dout <= -'sd2263; // 515
        'h204: dout <= -'sd740; // 516
        'h205: dout <=  'sd2033; // 517
        'h206: dout <=  'sd1299; // 518
        'h207: dout <= -'sd2123; // 519
        'h208: dout <= -'sd2043; // 520
        'h209: dout <= -'sd311; // 521
        'h20a: dout <= -'sd162; // 522
        'h20b: dout <= -'sd603; // 523
        'h20c: dout <= -'sd879; // 524
        'h20d: dout <=  'sd37; // 525
        'h20e: dout <= -'sd1080; // 526
        'h20f: dout <=  'sd2147; // 527
        'h210: dout <= -'sd653; // 528
        'h211: dout <= -'sd57; // 529
        'h212: dout <=  'sd253; // 530
        'h213: dout <= -'sd240; // 531
        'h214: dout <=  'sd1361; // 532
        'h215: dout <= -'sd919; // 533
        'h216: dout <=  'sd2172; // 534
        'h217: dout <=  'sd629; // 535
        'h218: dout <=  'sd1725; // 536
        'h219: dout <=  'sd1145; // 537
        'h21a: dout <= -'sd1298; // 538
        'h21b: dout <= -'sd584; // 539
        'h21c: dout <=  'sd844; // 540
        'h21d: dout <= -'sd618; // 541
        'h21e: dout <=  'sd31; // 542
        'h21f: dout <= -'sd1410; // 543
        'h220: dout <= -'sd2098; // 544
        'h221: dout <= -'sd1328; // 545
        'h222: dout <= -'sd2187; // 546
        'h223: dout <=  'sd2171; // 547
        'h224: dout <=  'sd133; // 548
        'h225: dout <= -'sd1177; // 549
        'h226: dout <= -'sd1680; // 550
        'h227: dout <=  'sd1804; // 551
        'h228: dout <=  'sd766; // 552
        'h229: dout <=  'sd254; // 553
        'h22a: dout <=  'sd1286; // 554
        'h22b: dout <=  'sd1825; // 555
        'h22c: dout <=  'sd628; // 556
        'h22d: dout <=  'sd2033; // 557
        'h22e: dout <=  'sd356; // 558
        'h22f: dout <= -'sd2289; // 559
        'h230: dout <= -'sd1281; // 560
        'h231: dout <=  'sd1328; // 561
        'h232: dout <=  'sd1387; // 562
        'h233: dout <=  'sd573; // 563
        'h234: dout <=  'sd201; // 564
        'h235: dout <=  'sd2122; // 565
        'h236: dout <=  'sd976; // 566
        'h237: dout <=  'sd485; // 567
        'h238: dout <=  'sd1737; // 568
        'h239: dout <= -'sd1369; // 569
        'h23a: dout <=  'sd797; // 570
        'h23b: dout <=  'sd837; // 571
        'h23c: dout <= -'sd625; // 572
        'h23d: dout <=  'sd2267; // 573
        'h23e: dout <= -'sd2264; // 574
        'h23f: dout <= -'sd21; // 575
        'h240: dout <=  'sd1890; // 576
        'h241: dout <= -'sd666; // 577
        'h242: dout <=  'sd1486; // 578
        'h243: dout <=  'sd1939; // 579
        'h244: dout <=  'sd1055; // 580
        'h245: dout <=  'sd206; // 581
        'h246: dout <= -'sd900; // 582
        'h247: dout <=  'sd1386; // 583
        'h248: dout <=  'sd2054; // 584
        'h249: dout <= -'sd679; // 585
        'h24a: dout <=  'sd649; // 586
        'h24b: dout <=  'sd2015; // 587
        'h24c: dout <= -'sd2267; // 588
        'h24d: dout <=  'sd893; // 589
        'h24e: dout <=  'sd1193; // 590
        'h24f: dout <=  'sd1024; // 591
        'h250: dout <=  'sd457; // 592
        'h251: dout <= -'sd1741; // 593
        'h252: dout <=  'sd1741; // 594
        'h253: dout <= -'sd267; // 595
        'h254: dout <=  'sd87; // 596
        'h255: dout <= -'sd2125; // 597
        'h256: dout <=  'sd1039; // 598
        'h257: dout <= -'sd1017; // 599
        'h258: dout <=  'sd959; // 600
        'h259: dout <= -'sd82; // 601
        'h25a: dout <= -'sd836; // 602
        'h25b: dout <= -'sd1694; // 603
        'h25c: dout <= -'sd2213; // 604
        'h25d: dout <=  'sd567; // 605
        'h25e: dout <= -'sd128; // 606
        'h25f: dout <=  'sd1073; // 607
        'h260: dout <=  'sd2163; // 608
        'h261: dout <=  'sd192; // 609
        'h262: dout <= -'sd1050; // 610
        'h263: dout <=  'sd1490; // 611
        'h264: dout <= -'sd171; // 612
        'h265: dout <=  'sd1674; // 613
        'h266: dout <= -'sd906; // 614
        'h267: dout <=  'sd1531; // 615
        'h268: dout <=  'sd1885; // 616
        'h269: dout <= -'sd1924; // 617
        'h26a: dout <= -'sd77; // 618
        'h26b: dout <=  'sd1885; // 619
        'h26c: dout <= -'sd1488; // 620
        'h26d: dout <=  'sd1166; // 621
        'h26e: dout <= -'sd1724; // 622
        'h26f: dout <=  'sd614; // 623
        'h270: dout <= -'sd1747; // 624
        'h271: dout <=  'sd1329; // 625
        'h272: dout <= -'sd2134; // 626
        'h273: dout <= -'sd951; // 627
        'h274: dout <=  'sd1859; // 628
        'h275: dout <= -'sd971; // 629
        'h276: dout <= -'sd1533; // 630
        'h277: dout <=  'sd997; // 631
        'h278: dout <= -'sd36; // 632
        'h279: dout <=  'sd198; // 633
        'h27a: dout <= -'sd584; // 634
        'h27b: dout <=  'sd2031; // 635
        'h27c: dout <= -'sd594; // 636
        'h27d: dout <= -'sd352; // 637
        'h27e: dout <=  'sd440; // 638
        'h27f: dout <= -'sd91; // 639
        'h280: dout <= -'sd1734; // 640
        'h281: dout <= -'sd1682; // 641
        'h282: dout <=  'sd1991; // 642
        'h283: dout <=  'sd721; // 643
        'h284: dout <=  'sd1538; // 644
        'h285: dout <=  'sd1895; // 645
        'h286: dout <=  'sd2273; // 646
        'h287: dout <= -'sd1888; // 647
        'h288: dout <= -'sd915; // 648
        'h289: dout <=  'sd137; // 649
        'h28a: dout <=  'sd2261; // 650
        'h28b: dout <= -'sd86; // 651
        'h28c: dout <=  'sd620; // 652
        'h28d: dout <= -'sd394; // 653
        'h28e: dout <=  'sd920; // 654
        'h28f: dout <=  'sd979; // 655
        'h290: dout <= -'sd884; // 656
        'h291: dout <=  'sd1666; // 657
        'h292: dout <= -'sd169; // 658
        'h293: dout <=  'sd405; // 659
        'h294: dout <= -'sd474; // 660
        'h295: dout <= -'sd176; // 661
        'h296: dout <= -'sd295; // 662
        'h297: dout <= -'sd2045; // 663
        'h298: dout <=  'sd1003; // 664
        'h299: dout <=  'sd298; // 665
        'h29a: dout <=  'sd1242; // 666
        'h29b: dout <= -'sd260; // 667
        'h29c: dout <= -'sd91; // 668
        'h29d: dout <= -'sd740; // 669
        'h29e: dout <= -'sd1701; // 670
        'h29f: dout <= -'sd939; // 671
        'h2a0: dout <=  'sd1338; // 672
        'h2a1: dout <= -'sd1082; // 673
        'h2a2: dout <= -'sd149; // 674
        'h2a3: dout <=  'sd1468; // 675
        'h2a4: dout <=  'sd2018; // 676
        'h2a5: dout <= -'sd964; // 677
        'h2a6: dout <= -'sd1160; // 678
        'h2a7: dout <= -'sd1164; // 679
        'h2a8: dout <=  'sd1315; // 680
        'h2a9: dout <=  'sd663; // 681
        'h2aa: dout <=  'sd242; // 682
        'h2ab: dout <=  'sd987; // 683
        'h2ac: dout <= -'sd325; // 684
        'h2ad: dout <= -'sd1347; // 685
        'h2ae: dout <= -'sd606; // 686
        'h2af: dout <=  'sd207; // 687
        'h2b0: dout <= -'sd1737; // 688
        'h2b1: dout <= -'sd1424; // 689
        'h2b2: dout <= -'sd431; // 690
        'h2b3: dout <=  'sd957; // 691
        'h2b4: dout <=  'sd337; // 692
        'h2b5: dout <=  'sd1738; // 693
        'h2b6: dout <= -'sd1477; // 694
        'h2b7: dout <= -'sd766; // 695
        'h2b8: dout <= -'sd1927; // 696
        'h2b9: dout <= -'sd1842; // 697
        'h2ba: dout <= -'sd2105; // 698
        'h2bb: dout <= -'sd521; // 699
        'h2bc: dout <= -'sd2011; // 700
        'h2bd: dout <=  'sd1755; // 701
        'h2be: dout <=  'sd2034; // 702
        'h2bf: dout <=  'sd1328; // 703
        'h2c0: dout <=  'sd510; // 704
        'h2c1: dout <= -'sd46; // 705
        'h2c2: dout <= -'sd1328; // 706
        'h2c3: dout <= -'sd881; // 707
        'h2c4: dout <= -'sd1515; // 708
        'h2c5: dout <= -'sd476; // 709
        'h2c6: dout <=  'sd979; // 710
        'h2c7: dout <= -'sd385; // 711
        'h2c8: dout <=  'sd1760; // 712
        'h2c9: dout <=  'sd1389; // 713
        'h2ca: dout <=  'sd800; // 714
        'h2cb: dout <= -'sd914; // 715
        'h2cc: dout <= -'sd397; // 716
        'h2cd: dout <= -'sd364; // 717
        'h2ce: dout <=  'sd28; // 718
        'h2cf: dout <=  'sd1494; // 719
        'h2d0: dout <=  'sd2186; // 720
        'h2d1: dout <=  'sd896; // 721
        'h2d2: dout <= -'sd560; // 722
        'h2d3: dout <=  'sd1405; // 723
        'h2d4: dout <= -'sd183; // 724
        'h2d5: dout <=  'sd409; // 725
        'h2d6: dout <=  'sd1770; // 726
        'h2d7: dout <= -'sd1387; // 727
        'h2d8: dout <= -'sd544; // 728
        'h2d9: dout <= -'sd1650; // 729
        'h2da: dout <= -'sd1917; // 730
        'h2db: dout <= -'sd2169; // 731
        'h2dc: dout <= -'sd2253; // 732
        'h2dd: dout <=  'sd1640; // 733
        'h2de: dout <=  'sd322; // 734
        'h2df: dout <=  'sd843; // 735
        'h2e0: dout <=  'sd57; // 736
        'h2e1: dout <= -'sd691; // 737
        'h2e2: dout <=  'sd981; // 738
        'h2e3: dout <= -'sd984; // 739
        'h2e4: dout <= -'sd1048; // 740
        'h2e5: dout <= -'sd2046; // 741
        'h2e6: dout <= -'sd2171; // 742
        'h2e7: dout <=  'sd877; // 743
        'h2e8: dout <= -'sd1106; // 744
        'h2e9: dout <=  'sd2149; // 745
        'h2ea: dout <= -'sd1828; // 746
        'h2eb: dout <=  'sd813; // 747
        'h2ec: dout <= -'sd213; // 748
        'h2ed: dout <= -'sd1231; // 749
        'h2ee: dout <= -'sd1644; // 750
        'h2ef: dout <=  'sd1496; // 751
        'h2f0: dout <=  'sd190; // 752
        'h2f1: dout <= -'sd2177; // 753
        'h2f2: dout <= -'sd2005; // 754
        'h2f3: dout <=  'sd2103; // 755
        'h2f4: dout <= -'sd1797; // 756
        'h2f5: dout <=  'sd2005; // 757
        'h2f6: dout <= -'sd1239; // 758
        'h2f7: dout <= -'sd1945; // 759
        'h2f8: dout <= -'sd54; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module g_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [12:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd1333; // 0
        'h001: dout <=  'sd1248; // 1
        'h002: dout <= -'sd1550; // 2
        'h003: dout <= -'sd738; // 3
        'h004: dout <= -'sd2069; // 4
        'h005: dout <=  'sd1798; // 5
        'h006: dout <= -'sd1228; // 6
        'h007: dout <= -'sd8; // 7
        'h008: dout <= -'sd723; // 8
        'h009: dout <=  'sd1371; // 9
        'h00a: dout <=  'sd897; // 10
        'h00b: dout <=  'sd406; // 11
        'h00c: dout <= -'sd100; // 12
        'h00d: dout <= -'sd167; // 13
        'h00e: dout <= -'sd304; // 14
        'h00f: dout <= -'sd285; // 15
        'h010: dout <= -'sd1802; // 16
        'h011: dout <= -'sd860; // 17
        'h012: dout <=  'sd569; // 18
        'h013: dout <=  'sd1215; // 19
        'h014: dout <=  'sd2294; // 20
        'h015: dout <=  'sd1982; // 21
        'h016: dout <= -'sd1797; // 22
        'h017: dout <=  'sd598; // 23
        'h018: dout <=  'sd2185; // 24
        'h019: dout <=  'sd1085; // 25
        'h01a: dout <=  'sd2113; // 26
        'h01b: dout <= -'sd662; // 27
        'h01c: dout <=  'sd2099; // 28
        'h01d: dout <=  'sd1179; // 29
        'h01e: dout <= -'sd1721; // 30
        'h01f: dout <= -'sd107; // 31
        'h020: dout <= -'sd1703; // 32
        'h021: dout <= -'sd235; // 33
        'h022: dout <= -'sd841; // 34
        'h023: dout <= -'sd1504; // 35
        'h024: dout <= -'sd1058; // 36
        'h025: dout <= -'sd1815; // 37
        'h026: dout <= -'sd630; // 38
        'h027: dout <=  'sd1212; // 39
        'h028: dout <= -'sd1928; // 40
        'h029: dout <= -'sd1863; // 41
        'h02a: dout <= -'sd1548; // 42
        'h02b: dout <=  'sd1906; // 43
        'h02c: dout <=  'sd1548; // 44
        'h02d: dout <=  'sd1810; // 45
        'h02e: dout <=  'sd738; // 46
        'h02f: dout <= -'sd1482; // 47
        'h030: dout <=  'sd266; // 48
        'h031: dout <= -'sd1967; // 49
        'h032: dout <= -'sd1258; // 50
        'h033: dout <=  'sd2058; // 51
        'h034: dout <= -'sd2024; // 52
        'h035: dout <=  'sd1336; // 53
        'h036: dout <= -'sd1245; // 54
        'h037: dout <=  'sd942; // 55
        'h038: dout <=  'sd1359; // 56
        'h039: dout <= -'sd2094; // 57
        'h03a: dout <=  'sd2001; // 58
        'h03b: dout <= -'sd84; // 59
        'h03c: dout <= -'sd1555; // 60
        'h03d: dout <= -'sd247; // 61
        'h03e: dout <=  'sd370; // 62
        'h03f: dout <= -'sd1593; // 63
        'h040: dout <=  'sd177; // 64
        'h041: dout <= -'sd2015; // 65
        'h042: dout <=  'sd852; // 66
        'h043: dout <= -'sd1819; // 67
        'h044: dout <= -'sd157; // 68
        'h045: dout <=  'sd270; // 69
        'h046: dout <= -'sd1230; // 70
        'h047: dout <= -'sd163; // 71
        'h048: dout <=  'sd819; // 72
        'h049: dout <= -'sd1336; // 73
        'h04a: dout <=  'sd193; // 74
        'h04b: dout <= -'sd1525; // 75
        'h04c: dout <=  'sd1185; // 76
        'h04d: dout <= -'sd285; // 77
        'h04e: dout <=  'sd1823; // 78
        'h04f: dout <=  'sd2269; // 79
        'h050: dout <= -'sd613; // 80
        'h051: dout <=  'sd409; // 81
        'h052: dout <=  'sd479; // 82
        'h053: dout <=  'sd1877; // 83
        'h054: dout <=  'sd908; // 84
        'h055: dout <=  'sd1646; // 85
        'h056: dout <= -'sd1438; // 86
        'h057: dout <= -'sd1233; // 87
        'h058: dout <=  'sd1380; // 88
        'h059: dout <=  'sd1995; // 89
        'h05a: dout <=  'sd2281; // 90
        'h05b: dout <=  'sd1965; // 91
        'h05c: dout <=  'sd2092; // 92
        'h05d: dout <= -'sd2048; // 93
        'h05e: dout <=  'sd91; // 94
        'h05f: dout <= -'sd1009; // 95
        'h060: dout <= -'sd657; // 96
        'h061: dout <=  'sd738; // 97
        'h062: dout <=  'sd893; // 98
        'h063: dout <=  'sd1973; // 99
        'h064: dout <=  'sd361; // 100
        'h065: dout <= -'sd1498; // 101
        'h066: dout <=  'sd1059; // 102
        'h067: dout <=  'sd534; // 103
        'h068: dout <= -'sd1260; // 104
        'h069: dout <= -'sd1764; // 105
        'h06a: dout <= -'sd1939; // 106
        'h06b: dout <=  'sd166; // 107
        'h06c: dout <=  'sd2076; // 108
        'h06d: dout <=  'sd274; // 109
        'h06e: dout <=  'sd1125; // 110
        'h06f: dout <=  'sd148; // 111
        'h070: dout <=  'sd316; // 112
        'h071: dout <=  'sd593; // 113
        'h072: dout <= -'sd62; // 114
        'h073: dout <=  'sd369; // 115
        'h074: dout <=  'sd1965; // 116
        'h075: dout <=  'sd1809; // 117
        'h076: dout <= -'sd2225; // 118
        'h077: dout <=  'sd2015; // 119
        'h078: dout <= -'sd1297; // 120
        'h079: dout <= -'sd1077; // 121
        'h07a: dout <=  'sd302; // 122
        'h07b: dout <=  'sd372; // 123
        'h07c: dout <=  'sd388; // 124
        'h07d: dout <= -'sd1732; // 125
        'h07e: dout <=  'sd1406; // 126
        'h07f: dout <= -'sd5; // 127
        'h080: dout <=  'sd1634; // 128
        'h081: dout <=  'sd1425; // 129
        'h082: dout <=  'sd688; // 130
        'h083: dout <=  'sd822; // 131
        'h084: dout <= -'sd1655; // 132
        'h085: dout <= -'sd1836; // 133
        'h086: dout <= -'sd1193; // 134
        'h087: dout <= -'sd1896; // 135
        'h088: dout <=  'sd1995; // 136
        'h089: dout <=  'sd1736; // 137
        'h08a: dout <= -'sd232; // 138
        'h08b: dout <= -'sd285; // 139
        'h08c: dout <=  'sd479; // 140
        'h08d: dout <=  'sd667; // 141
        'h08e: dout <=  'sd737; // 142
        'h08f: dout <=  'sd1002; // 143
        'h090: dout <=  'sd223; // 144
        'h091: dout <=  'sd1510; // 145
        'h092: dout <=  'sd493; // 146
        'h093: dout <=  'sd2064; // 147
        'h094: dout <=  'sd1862; // 148
        'h095: dout <= -'sd921; // 149
        'h096: dout <= -'sd2057; // 150
        'h097: dout <= -'sd1080; // 151
        'h098: dout <= -'sd246; // 152
        'h099: dout <= -'sd484; // 153
        'h09a: dout <= -'sd1203; // 154
        'h09b: dout <= -'sd1372; // 155
        'h09c: dout <= -'sd783; // 156
        'h09d: dout <=  'sd1072; // 157
        'h09e: dout <= -'sd1885; // 158
        'h09f: dout <= -'sd1483; // 159
        'h0a0: dout <=  'sd2175; // 160
        'h0a1: dout <= -'sd119; // 161
        'h0a2: dout <= -'sd1419; // 162
        'h0a3: dout <= -'sd622; // 163
        'h0a4: dout <= -'sd152; // 164
        'h0a5: dout <= -'sd1748; // 165
        'h0a6: dout <=  'sd2017; // 166
        'h0a7: dout <= -'sd1652; // 167
        'h0a8: dout <= -'sd1699; // 168
        'h0a9: dout <= -'sd515; // 169
        'h0aa: dout <= -'sd875; // 170
        'h0ab: dout <=  'sd1895; // 171
        'h0ac: dout <=  'sd1244; // 172
        'h0ad: dout <= -'sd2117; // 173
        'h0ae: dout <=  'sd720; // 174
        'h0af: dout <=  'sd1691; // 175
        'h0b0: dout <=  'sd29; // 176
        'h0b1: dout <= -'sd494; // 177
        'h0b2: dout <= -'sd654; // 178
        'h0b3: dout <=  'sd1748; // 179
        'h0b4: dout <= -'sd369; // 180
        'h0b5: dout <=  'sd1190; // 181
        'h0b6: dout <=  'sd1409; // 182
        'h0b7: dout <=  'sd712; // 183
        'h0b8: dout <=  'sd2165; // 184
        'h0b9: dout <= -'sd749; // 185
        'h0ba: dout <=  'sd1654; // 186
        'h0bb: dout <= -'sd1700; // 187
        'h0bc: dout <= -'sd194; // 188
        'h0bd: dout <=  'sd1041; // 189
        'h0be: dout <= -'sd646; // 190
        'h0bf: dout <= -'sd2228; // 191
        'h0c0: dout <=  'sd2063; // 192
        'h0c1: dout <=  'sd823; // 193
        'h0c2: dout <=  'sd1918; // 194
        'h0c3: dout <=  'sd1695; // 195
        'h0c4: dout <= -'sd1670; // 196
        'h0c5: dout <=  'sd1012; // 197
        'h0c6: dout <=  'sd1883; // 198
        'h0c7: dout <=  'sd1191; // 199
        'h0c8: dout <= -'sd1967; // 200
        'h0c9: dout <=  'sd587; // 201
        'h0ca: dout <=  'sd1460; // 202
        'h0cb: dout <= -'sd2243; // 203
        'h0cc: dout <= -'sd741; // 204
        'h0cd: dout <=  'sd157; // 205
        'h0ce: dout <= -'sd2250; // 206
        'h0cf: dout <=  'sd2135; // 207
        'h0d0: dout <= -'sd1312; // 208
        'h0d1: dout <=  'sd184; // 209
        'h0d2: dout <=  'sd1903; // 210
        'h0d3: dout <=  'sd290; // 211
        'h0d4: dout <=  'sd2153; // 212
        'h0d5: dout <=  'sd2221; // 213
        'h0d6: dout <=  'sd19; // 214
        'h0d7: dout <=  'sd2010; // 215
        'h0d8: dout <=  'sd1075; // 216
        'h0d9: dout <=  'sd2145; // 217
        'h0da: dout <=  'sd1947; // 218
        'h0db: dout <=  'sd1049; // 219
        'h0dc: dout <=  'sd226; // 220
        'h0dd: dout <=  'sd1412; // 221
        'h0de: dout <=  'sd178; // 222
        'h0df: dout <= -'sd1223; // 223
        'h0e0: dout <=  'sd1852; // 224
        'h0e1: dout <=  'sd1343; // 225
        'h0e2: dout <= -'sd1146; // 226
        'h0e3: dout <=  'sd2210; // 227
        'h0e4: dout <= -'sd960; // 228
        'h0e5: dout <= -'sd225; // 229
        'h0e6: dout <= -'sd2217; // 230
        'h0e7: dout <=  'sd1179; // 231
        'h0e8: dout <= -'sd1999; // 232
        'h0e9: dout <=  'sd722; // 233
        'h0ea: dout <=  'sd1152; // 234
        'h0eb: dout <=  'sd999; // 235
        'h0ec: dout <=  'sd11; // 236
        'h0ed: dout <= -'sd2145; // 237
        'h0ee: dout <= -'sd1554; // 238
        'h0ef: dout <= -'sd1558; // 239
        'h0f0: dout <= -'sd2256; // 240
        'h0f1: dout <=  'sd845; // 241
        'h0f2: dout <= -'sd93; // 242
        'h0f3: dout <=  'sd1509; // 243
        'h0f4: dout <= -'sd68; // 244
        'h0f5: dout <=  'sd757; // 245
        'h0f6: dout <=  'sd1648; // 246
        'h0f7: dout <=  'sd461; // 247
        'h0f8: dout <=  'sd887; // 248
        'h0f9: dout <=  'sd1441; // 249
        'h0fa: dout <= -'sd1341; // 250
        'h0fb: dout <=  'sd1667; // 251
        'h0fc: dout <=  'sd609; // 252
        'h0fd: dout <= -'sd1110; // 253
        'h0fe: dout <=  'sd1106; // 254
        'h0ff: dout <= -'sd1081; // 255
        'h100: dout <= -'sd2147; // 256
        'h101: dout <= -'sd886; // 257
        'h102: dout <= -'sd164; // 258
        'h103: dout <=  'sd717; // 259
        'h104: dout <= -'sd1254; // 260
        'h105: dout <=  'sd57; // 261
        'h106: dout <=  'sd1087; // 262
        'h107: dout <= -'sd183; // 263
        'h108: dout <=  'sd1913; // 264
        'h109: dout <=  'sd58; // 265
        'h10a: dout <=  'sd1151; // 266
        'h10b: dout <= -'sd54; // 267
        'h10c: dout <=  'sd1256; // 268
        'h10d: dout <=  'sd456; // 269
        'h10e: dout <=  'sd1684; // 270
        'h10f: dout <= -'sd530; // 271
        'h110: dout <=  'sd1730; // 272
        'h111: dout <=  'sd997; // 273
        'h112: dout <=  'sd1187; // 274
        'h113: dout <= -'sd1547; // 275
        'h114: dout <= -'sd1768; // 276
        'h115: dout <= -'sd1235; // 277
        'h116: dout <= -'sd607; // 278
        'h117: dout <= -'sd1070; // 279
        'h118: dout <= -'sd418; // 280
        'h119: dout <= -'sd2081; // 281
        'h11a: dout <= -'sd1450; // 282
        'h11b: dout <= -'sd221; // 283
        'h11c: dout <= -'sd1020; // 284
        'h11d: dout <=  'sd1635; // 285
        'h11e: dout <= -'sd1485; // 286
        'h11f: dout <=  'sd974; // 287
        'h120: dout <= -'sd760; // 288
        'h121: dout <= -'sd2271; // 289
        'h122: dout <= -'sd1565; // 290
        'h123: dout <=  'sd1208; // 291
        'h124: dout <= -'sd1879; // 292
        'h125: dout <=  'sd2207; // 293
        'h126: dout <= -'sd507; // 294
        'h127: dout <=  'sd2083; // 295
        'h128: dout <=  'sd1161; // 296
        'h129: dout <=  'sd545; // 297
        'h12a: dout <= -'sd1910; // 298
        'h12b: dout <= -'sd1450; // 299
        'h12c: dout <=  'sd2233; // 300
        'h12d: dout <=  'sd1142; // 301
        'h12e: dout <= -'sd1324; // 302
        'h12f: dout <= -'sd122; // 303
        'h130: dout <= -'sd12; // 304
        'h131: dout <= -'sd829; // 305
        'h132: dout <=  'sd1634; // 306
        'h133: dout <= -'sd1905; // 307
        'h134: dout <= -'sd541; // 308
        'h135: dout <= -'sd1581; // 309
        'h136: dout <=  'sd897; // 310
        'h137: dout <= -'sd1281; // 311
        'h138: dout <=  'sd1369; // 312
        'h139: dout <=  'sd115; // 313
        'h13a: dout <=  'sd1865; // 314
        'h13b: dout <=  'sd1784; // 315
        'h13c: dout <=  'sd925; // 316
        'h13d: dout <= -'sd1344; // 317
        'h13e: dout <=  'sd1630; // 318
        'h13f: dout <= -'sd1429; // 319
        'h140: dout <= -'sd1074; // 320
        'h141: dout <=  'sd870; // 321
        'h142: dout <= -'sd647; // 322
        'h143: dout <= -'sd926; // 323
        'h144: dout <=  'sd1970; // 324
        'h145: dout <= -'sd185; // 325
        'h146: dout <=  'sd1117; // 326
        'h147: dout <=  'sd2101; // 327
        'h148: dout <=  'sd69; // 328
        'h149: dout <=  'sd1739; // 329
        'h14a: dout <=  'sd2167; // 330
        'h14b: dout <= -'sd537; // 331
        'h14c: dout <=  'sd466; // 332
        'h14d: dout <=  'sd1686; // 333
        'h14e: dout <= -'sd1453; // 334
        'h14f: dout <= -'sd2225; // 335
        'h150: dout <=  'sd546; // 336
        'h151: dout <= -'sd104; // 337
        'h152: dout <= -'sd1833; // 338
        'h153: dout <=  'sd2133; // 339
        'h154: dout <=  'sd1311; // 340
        'h155: dout <=  'sd161; // 341
        'h156: dout <= -'sd1470; // 342
        'h157: dout <= -'sd423; // 343
        'h158: dout <=  'sd1866; // 344
        'h159: dout <= -'sd46; // 345
        'h15a: dout <= -'sd81; // 346
        'h15b: dout <= -'sd277; // 347
        'h15c: dout <=  'sd1077; // 348
        'h15d: dout <= -'sd1080; // 349
        'h15e: dout <= -'sd1229; // 350
        'h15f: dout <= -'sd196; // 351
        'h160: dout <= -'sd696; // 352
        'h161: dout <=  'sd1045; // 353
        'h162: dout <= -'sd1817; // 354
        'h163: dout <=  'sd2069; // 355
        'h164: dout <=  'sd1877; // 356
        'h165: dout <= -'sd1076; // 357
        'h166: dout <=  'sd1094; // 358
        'h167: dout <= -'sd82; // 359
        'h168: dout <= -'sd3; // 360
        'h169: dout <=  'sd1638; // 361
        'h16a: dout <=  'sd210; // 362
        'h16b: dout <= -'sd108; // 363
        'h16c: dout <=  'sd1729; // 364
        'h16d: dout <= -'sd539; // 365
        'h16e: dout <=  'sd1790; // 366
        'h16f: dout <=  'sd717; // 367
        'h170: dout <=  'sd1559; // 368
        'h171: dout <= -'sd316; // 369
        'h172: dout <=  'sd477; // 370
        'h173: dout <= -'sd852; // 371
        'h174: dout <= -'sd811; // 372
        'h175: dout <=  'sd1400; // 373
        'h176: dout <=  'sd2085; // 374
        'h177: dout <= -'sd1071; // 375
        'h178: dout <= -'sd1819; // 376
        'h179: dout <=  'sd1833; // 377
        'h17a: dout <=  'sd375; // 378
        'h17b: dout <=  'sd2034; // 379
        'h17c: dout <= -'sd1189; // 380
        'h17d: dout <= -'sd549; // 381
        'h17e: dout <=  'sd288; // 382
        'h17f: dout <=  'sd1749; // 383
        'h180: dout <=  'sd1640; // 384
        'h181: dout <=  'sd408; // 385
        'h182: dout <= -'sd1326; // 386
        'h183: dout <= -'sd1248; // 387
        'h184: dout <= -'sd1148; // 388
        'h185: dout <= -'sd195; // 389
        'h186: dout <= -'sd452; // 390
        'h187: dout <= -'sd1574; // 391
        'h188: dout <=  'sd2119; // 392
        'h189: dout <= -'sd1886; // 393
        'h18a: dout <= -'sd886; // 394
        'h18b: dout <= -'sd1344; // 395
        'h18c: dout <= -'sd442; // 396
        'h18d: dout <= -'sd662; // 397
        'h18e: dout <=  'sd1825; // 398
        'h18f: dout <=  'sd227; // 399
        'h190: dout <=  'sd1164; // 400
        'h191: dout <=  'sd389; // 401
        'h192: dout <= -'sd2261; // 402
        'h193: dout <= -'sd2131; // 403
        'h194: dout <=  'sd206; // 404
        'h195: dout <= -'sd491; // 405
        'h196: dout <= -'sd1603; // 406
        'h197: dout <= -'sd456; // 407
        'h198: dout <=  'sd0; // 408
        'h199: dout <=  'sd499; // 409
        'h19a: dout <= -'sd91; // 410
        'h19b: dout <=  'sd1951; // 411
        'h19c: dout <=  'sd812; // 412
        'h19d: dout <= -'sd2106; // 413
        'h19e: dout <= -'sd1299; // 414
        'h19f: dout <=  'sd407; // 415
        'h1a0: dout <=  'sd547; // 416
        'h1a1: dout <= -'sd1153; // 417
        'h1a2: dout <= -'sd1367; // 418
        'h1a3: dout <= -'sd241; // 419
        'h1a4: dout <= -'sd1122; // 420
        'h1a5: dout <= -'sd1959; // 421
        'h1a6: dout <=  'sd547; // 422
        'h1a7: dout <= -'sd1662; // 423
        'h1a8: dout <= -'sd1543; // 424
        'h1a9: dout <= -'sd1450; // 425
        'h1aa: dout <=  'sd162; // 426
        'h1ab: dout <=  'sd302; // 427
        'h1ac: dout <= -'sd256; // 428
        'h1ad: dout <= -'sd89; // 429
        'h1ae: dout <=  'sd2043; // 430
        'h1af: dout <= -'sd1888; // 431
        'h1b0: dout <=  'sd668; // 432
        'h1b1: dout <= -'sd2040; // 433
        'h1b2: dout <= -'sd1654; // 434
        'h1b3: dout <= -'sd1157; // 435
        'h1b4: dout <=  'sd976; // 436
        'h1b5: dout <=  'sd752; // 437
        'h1b6: dout <= -'sd313; // 438
        'h1b7: dout <= -'sd1527; // 439
        'h1b8: dout <=  'sd398; // 440
        'h1b9: dout <= -'sd54; // 441
        'h1ba: dout <= -'sd2230; // 442
        'h1bb: dout <=  'sd1925; // 443
        'h1bc: dout <=  'sd341; // 444
        'h1bd: dout <= -'sd1376; // 445
        'h1be: dout <=  'sd591; // 446
        'h1bf: dout <= -'sd1264; // 447
        'h1c0: dout <= -'sd75; // 448
        'h1c1: dout <=  'sd1024; // 449
        'h1c2: dout <= -'sd1549; // 450
        'h1c3: dout <=  'sd2028; // 451
        'h1c4: dout <=  'sd1600; // 452
        'h1c5: dout <=  'sd1135; // 453
        'h1c6: dout <=  'sd2093; // 454
        'h1c7: dout <=  'sd930; // 455
        'h1c8: dout <=  'sd171; // 456
        'h1c9: dout <= -'sd498; // 457
        'h1ca: dout <=  'sd184; // 458
        'h1cb: dout <=  'sd2203; // 459
        'h1cc: dout <= -'sd1205; // 460
        'h1cd: dout <= -'sd1854; // 461
        'h1ce: dout <=  'sd1870; // 462
        'h1cf: dout <= -'sd1395; // 463
        'h1d0: dout <= -'sd861; // 464
        'h1d1: dout <= -'sd325; // 465
        'h1d2: dout <= -'sd534; // 466
        'h1d3: dout <=  'sd1265; // 467
        'h1d4: dout <= -'sd47; // 468
        'h1d5: dout <=  'sd2177; // 469
        'h1d6: dout <= -'sd2132; // 470
        'h1d7: dout <= -'sd244; // 471
        'h1d8: dout <=  'sd2119; // 472
        'h1d9: dout <= -'sd76; // 473
        'h1da: dout <=  'sd2047; // 474
        'h1db: dout <= -'sd151; // 475
        'h1dc: dout <=  'sd1581; // 476
        'h1dd: dout <= -'sd1263; // 477
        'h1de: dout <=  'sd1008; // 478
        'h1df: dout <= -'sd1446; // 479
        'h1e0: dout <=  'sd764; // 480
        'h1e1: dout <= -'sd1730; // 481
        'h1e2: dout <=  'sd2163; // 482
        'h1e3: dout <=  'sd679; // 483
        'h1e4: dout <=  'sd2167; // 484
        'h1e5: dout <=  'sd2255; // 485
        'h1e6: dout <=  'sd1861; // 486
        'h1e7: dout <= -'sd2046; // 487
        'h1e8: dout <=  'sd229; // 488
        'h1e9: dout <=  'sd1354; // 489
        'h1ea: dout <= -'sd1212; // 490
        'h1eb: dout <= -'sd1019; // 491
        'h1ec: dout <= -'sd1686; // 492
        'h1ed: dout <= -'sd1133; // 493
        'h1ee: dout <= -'sd524; // 494
        'h1ef: dout <=  'sd1670; // 495
        'h1f0: dout <=  'sd453; // 496
        'h1f1: dout <=  'sd695; // 497
        'h1f2: dout <=  'sd99; // 498
        'h1f3: dout <= -'sd987; // 499
        'h1f4: dout <= -'sd1021; // 500
        'h1f5: dout <=  'sd832; // 501
        'h1f6: dout <=  'sd1307; // 502
        'h1f7: dout <=  'sd1028; // 503
        'h1f8: dout <= -'sd1330; // 504
        'h1f9: dout <= -'sd1106; // 505
        'h1fa: dout <= -'sd86; // 506
        'h1fb: dout <=  'sd124; // 507
        'h1fc: dout <= -'sd2228; // 508
        'h1fd: dout <=  'sd2106; // 509
        'h1fe: dout <= -'sd2216; // 510
        'h1ff: dout <= -'sd1209; // 511
        'h200: dout <=  'sd813; // 512
        'h201: dout <= -'sd1467; // 513
        'h202: dout <=  'sd1469; // 514
        'h203: dout <= -'sd2047; // 515
        'h204: dout <=  'sd1243; // 516
        'h205: dout <=  'sd1164; // 517
        'h206: dout <= -'sd34; // 518
        'h207: dout <=  'sd737; // 519
        'h208: dout <=  'sd1050; // 520
        'h209: dout <=  'sd1032; // 521
        'h20a: dout <=  'sd1489; // 522
        'h20b: dout <= -'sd1859; // 523
        'h20c: dout <= -'sd1483; // 524
        'h20d: dout <=  'sd1561; // 525
        'h20e: dout <= -'sd1989; // 526
        'h20f: dout <= -'sd2291; // 527
        'h210: dout <= -'sd1951; // 528
        'h211: dout <= -'sd1385; // 529
        'h212: dout <= -'sd1152; // 530
        'h213: dout <=  'sd2050; // 531
        'h214: dout <=  'sd1867; // 532
        'h215: dout <=  'sd623; // 533
        'h216: dout <=  'sd2219; // 534
        'h217: dout <= -'sd76; // 535
        'h218: dout <=  'sd624; // 536
        'h219: dout <=  'sd1587; // 537
        'h21a: dout <= -'sd287; // 538
        'h21b: dout <= -'sd331; // 539
        'h21c: dout <= -'sd1431; // 540
        'h21d: dout <=  'sd635; // 541
        'h21e: dout <= -'sd996; // 542
        'h21f: dout <= -'sd1342; // 543
        'h220: dout <= -'sd1963; // 544
        'h221: dout <=  'sd274; // 545
        'h222: dout <=  'sd1165; // 546
        'h223: dout <=  'sd541; // 547
        'h224: dout <= -'sd219; // 548
        'h225: dout <= -'sd1839; // 549
        'h226: dout <=  'sd1267; // 550
        'h227: dout <=  'sd1104; // 551
        'h228: dout <=  'sd787; // 552
        'h229: dout <=  'sd643; // 553
        'h22a: dout <=  'sd112; // 554
        'h22b: dout <=  'sd500; // 555
        'h22c: dout <=  'sd1317; // 556
        'h22d: dout <= -'sd345; // 557
        'h22e: dout <=  'sd1956; // 558
        'h22f: dout <= -'sd1113; // 559
        'h230: dout <= -'sd1836; // 560
        'h231: dout <=  'sd502; // 561
        'h232: dout <= -'sd1366; // 562
        'h233: dout <=  'sd1907; // 563
        'h234: dout <= -'sd885; // 564
        'h235: dout <=  'sd2153; // 565
        'h236: dout <=  'sd1698; // 566
        'h237: dout <=  'sd498; // 567
        'h238: dout <= -'sd1300; // 568
        'h239: dout <= -'sd2118; // 569
        'h23a: dout <=  'sd1639; // 570
        'h23b: dout <= -'sd582; // 571
        'h23c: dout <=  'sd844; // 572
        'h23d: dout <= -'sd864; // 573
        'h23e: dout <=  'sd959; // 574
        'h23f: dout <= -'sd429; // 575
        'h240: dout <= -'sd1479; // 576
        'h241: dout <= -'sd261; // 577
        'h242: dout <=  'sd454; // 578
        'h243: dout <=  'sd400; // 579
        'h244: dout <= -'sd287; // 580
        'h245: dout <=  'sd1484; // 581
        'h246: dout <=  'sd1564; // 582
        'h247: dout <=  'sd732; // 583
        'h248: dout <=  'sd1740; // 584
        'h249: dout <= -'sd708; // 585
        'h24a: dout <=  'sd1243; // 586
        'h24b: dout <=  'sd1314; // 587
        'h24c: dout <=  'sd972; // 588
        'h24d: dout <=  'sd2145; // 589
        'h24e: dout <= -'sd1309; // 590
        'h24f: dout <=  'sd1704; // 591
        'h250: dout <= -'sd113; // 592
        'h251: dout <= -'sd1270; // 593
        'h252: dout <= -'sd1068; // 594
        'h253: dout <= -'sd2198; // 595
        'h254: dout <=  'sd786; // 596
        'h255: dout <=  'sd1101; // 597
        'h256: dout <= -'sd1403; // 598
        'h257: dout <= -'sd2081; // 599
        'h258: dout <= -'sd1684; // 600
        'h259: dout <= -'sd797; // 601
        'h25a: dout <=  'sd1463; // 602
        'h25b: dout <=  'sd793; // 603
        'h25c: dout <=  'sd1817; // 604
        'h25d: dout <=  'sd68; // 605
        'h25e: dout <= -'sd1022; // 606
        'h25f: dout <= -'sd1032; // 607
        'h260: dout <=  'sd2002; // 608
        'h261: dout <= -'sd1429; // 609
        'h262: dout <= -'sd210; // 610
        'h263: dout <= -'sd2142; // 611
        'h264: dout <=  'sd1509; // 612
        'h265: dout <=  'sd953; // 613
        'h266: dout <= -'sd425; // 614
        'h267: dout <=  'sd2110; // 615
        'h268: dout <=  'sd906; // 616
        'h269: dout <= -'sd2252; // 617
        'h26a: dout <=  'sd2162; // 618
        'h26b: dout <= -'sd252; // 619
        'h26c: dout <=  'sd1169; // 620
        'h26d: dout <= -'sd994; // 621
        'h26e: dout <= -'sd829; // 622
        'h26f: dout <=  'sd510; // 623
        'h270: dout <= -'sd336; // 624
        'h271: dout <= -'sd1672; // 625
        'h272: dout <=  'sd2098; // 626
        'h273: dout <=  'sd2274; // 627
        'h274: dout <= -'sd977; // 628
        'h275: dout <= -'sd857; // 629
        'h276: dout <=  'sd782; // 630
        'h277: dout <= -'sd2119; // 631
        'h278: dout <=  'sd1908; // 632
        'h279: dout <= -'sd519; // 633
        'h27a: dout <=  'sd1206; // 634
        'h27b: dout <= -'sd365; // 635
        'h27c: dout <= -'sd1964; // 636
        'h27d: dout <=  'sd1929; // 637
        'h27e: dout <= -'sd737; // 638
        'h27f: dout <=  'sd1834; // 639
        'h280: dout <=  'sd2102; // 640
        'h281: dout <= -'sd1663; // 641
        'h282: dout <= -'sd265; // 642
        'h283: dout <=  'sd966; // 643
        'h284: dout <=  'sd1513; // 644
        'h285: dout <= -'sd1320; // 645
        'h286: dout <= -'sd1899; // 646
        'h287: dout <=  'sd875; // 647
        'h288: dout <= -'sd1561; // 648
        'h289: dout <=  'sd2292; // 649
        'h28a: dout <= -'sd1521; // 650
        'h28b: dout <=  'sd1628; // 651
        'h28c: dout <= -'sd1927; // 652
        'h28d: dout <=  'sd1952; // 653
        'h28e: dout <= -'sd336; // 654
        'h28f: dout <= -'sd2196; // 655
        'h290: dout <= -'sd2125; // 656
        'h291: dout <=  'sd260; // 657
        'h292: dout <=  'sd1525; // 658
        'h293: dout <= -'sd18; // 659
        'h294: dout <=  'sd1109; // 660
        'h295: dout <= -'sd930; // 661
        'h296: dout <= -'sd1204; // 662
        'h297: dout <=  'sd312; // 663
        'h298: dout <=  'sd2085; // 664
        'h299: dout <=  'sd1380; // 665
        'h29a: dout <=  'sd1814; // 666
        'h29b: dout <=  'sd1126; // 667
        'h29c: dout <=  'sd2241; // 668
        'h29d: dout <= -'sd922; // 669
        'h29e: dout <=  'sd944; // 670
        'h29f: dout <=  'sd892; // 671
        'h2a0: dout <= -'sd651; // 672
        'h2a1: dout <=  'sd1763; // 673
        'h2a2: dout <= -'sd15; // 674
        'h2a3: dout <=  'sd654; // 675
        'h2a4: dout <= -'sd1055; // 676
        'h2a5: dout <= -'sd170; // 677
        'h2a6: dout <= -'sd6; // 678
        'h2a7: dout <= -'sd861; // 679
        'h2a8: dout <= -'sd1610; // 680
        'h2a9: dout <=  'sd658; // 681
        'h2aa: dout <=  'sd458; // 682
        'h2ab: dout <= -'sd1126; // 683
        'h2ac: dout <= -'sd178; // 684
        'h2ad: dout <= -'sd206; // 685
        'h2ae: dout <= -'sd229; // 686
        'h2af: dout <=  'sd566; // 687
        'h2b0: dout <=  'sd852; // 688
        'h2b1: dout <= -'sd9; // 689
        'h2b2: dout <=  'sd1536; // 690
        'h2b3: dout <= -'sd2185; // 691
        'h2b4: dout <= -'sd1075; // 692
        'h2b5: dout <= -'sd1228; // 693
        'h2b6: dout <= -'sd225; // 694
        'h2b7: dout <= -'sd445; // 695
        'h2b8: dout <= -'sd686; // 696
        'h2b9: dout <= -'sd1718; // 697
        'h2ba: dout <=  'sd2108; // 698
        'h2bb: dout <= -'sd670; // 699
        'h2bc: dout <=  'sd2153; // 700
        'h2bd: dout <=  'sd1221; // 701
        'h2be: dout <= -'sd331; // 702
        'h2bf: dout <= -'sd1155; // 703
        'h2c0: dout <=  'sd2242; // 704
        'h2c1: dout <=  'sd1477; // 705
        'h2c2: dout <=  'sd910; // 706
        'h2c3: dout <= -'sd691; // 707
        'h2c4: dout <= -'sd1619; // 708
        'h2c5: dout <= -'sd1663; // 709
        'h2c6: dout <= -'sd1041; // 710
        'h2c7: dout <= -'sd1824; // 711
        'h2c8: dout <= -'sd2048; // 712
        'h2c9: dout <=  'sd1025; // 713
        'h2ca: dout <=  'sd839; // 714
        'h2cb: dout <=  'sd1123; // 715
        'h2cc: dout <= -'sd1169; // 716
        'h2cd: dout <= -'sd1237; // 717
        'h2ce: dout <=  'sd2116; // 718
        'h2cf: dout <=  'sd2180; // 719
        'h2d0: dout <= -'sd1688; // 720
        'h2d1: dout <= -'sd319; // 721
        'h2d2: dout <=  'sd831; // 722
        'h2d3: dout <= -'sd1153; // 723
        'h2d4: dout <=  'sd45; // 724
        'h2d5: dout <= -'sd637; // 725
        'h2d6: dout <=  'sd958; // 726
        'h2d7: dout <=  'sd628; // 727
        'h2d8: dout <= -'sd835; // 728
        'h2d9: dout <= -'sd451; // 729
        'h2da: dout <=  'sd144; // 730
        'h2db: dout <= -'sd1117; // 731
        'h2dc: dout <=  'sd553; // 732
        'h2dd: dout <=  'sd1736; // 733
        'h2de: dout <=  'sd2090; // 734
        'h2df: dout <=  'sd95; // 735
        'h2e0: dout <= -'sd1570; // 736
        'h2e1: dout <=  'sd1918; // 737
        'h2e2: dout <=  'sd153; // 738
        'h2e3: dout <= -'sd585; // 739
        'h2e4: dout <=  'sd1501; // 740
        'h2e5: dout <= -'sd2116; // 741
        'h2e6: dout <=  'sd83; // 742
        'h2e7: dout <= -'sd1451; // 743
        'h2e8: dout <=  'sd757; // 744
        'h2e9: dout <=  'sd1338; // 745
        'h2ea: dout <= -'sd207; // 746
        'h2eb: dout <= -'sd1818; // 747
        'h2ec: dout <= -'sd1869; // 748
        'h2ed: dout <=  'sd290; // 749
        'h2ee: dout <= -'sd986; // 750
        'h2ef: dout <= -'sd1211; // 751
        'h2f0: dout <= -'sd1449; // 752
        'h2f1: dout <= -'sd1374; // 753
        'h2f2: dout <=  'sd1270; // 754
        'h2f3: dout <= -'sd281; // 755
        'h2f4: dout <= -'sd593; // 756
        'h2f5: dout <=  'sd1835; // 757
        'h2f6: dout <=  'sd1864; // 758
        'h2f7: dout <=  'sd955; // 759
        'h2f8: dout <= -'sd1300; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module h_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [12:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd142; // 0
        'h001: dout <= -'sd1425; // 1
        'h002: dout <= -'sd1524; // 2
        'h003: dout <= -'sd531; // 3
        'h004: dout <= -'sd1673; // 4
        'h005: dout <=  'sd1850; // 5
        'h006: dout <= -'sd1616; // 6
        'h007: dout <=  'sd976; // 7
        'h008: dout <=  'sd2207; // 8
        'h009: dout <= -'sd464; // 9
        'h00a: dout <=  'sd1801; // 10
        'h00b: dout <=  'sd1495; // 11
        'h00c: dout <=  'sd2281; // 12
        'h00d: dout <= -'sd2073; // 13
        'h00e: dout <=  'sd1602; // 14
        'h00f: dout <= -'sd1021; // 15
        'h010: dout <= -'sd119; // 16
        'h011: dout <=  'sd430; // 17
        'h012: dout <=  'sd500; // 18
        'h013: dout <= -'sd136; // 19
        'h014: dout <=  'sd884; // 20
        'h015: dout <= -'sd1565; // 21
        'h016: dout <= -'sd2183; // 22
        'h017: dout <= -'sd2222; // 23
        'h018: dout <= -'sd27; // 24
        'h019: dout <=  'sd1039; // 25
        'h01a: dout <=  'sd2273; // 26
        'h01b: dout <= -'sd1990; // 27
        'h01c: dout <= -'sd1124; // 28
        'h01d: dout <= -'sd1092; // 29
        'h01e: dout <= -'sd1678; // 30
        'h01f: dout <= -'sd114; // 31
        'h020: dout <= -'sd965; // 32
        'h021: dout <= -'sd219; // 33
        'h022: dout <=  'sd1056; // 34
        'h023: dout <= -'sd676; // 35
        'h024: dout <= -'sd369; // 36
        'h025: dout <= -'sd194; // 37
        'h026: dout <=  'sd645; // 38
        'h027: dout <= -'sd1225; // 39
        'h028: dout <= -'sd1103; // 40
        'h029: dout <=  'sd1459; // 41
        'h02a: dout <= -'sd937; // 42
        'h02b: dout <= -'sd1079; // 43
        'h02c: dout <=  'sd2211; // 44
        'h02d: dout <=  'sd1659; // 45
        'h02e: dout <= -'sd70; // 46
        'h02f: dout <= -'sd978; // 47
        'h030: dout <=  'sd1262; // 48
        'h031: dout <= -'sd1098; // 49
        'h032: dout <=  'sd1529; // 50
        'h033: dout <=  'sd1455; // 51
        'h034: dout <= -'sd333; // 52
        'h035: dout <=  'sd1577; // 53
        'h036: dout <=  'sd2086; // 54
        'h037: dout <= -'sd1878; // 55
        'h038: dout <= -'sd1486; // 56
        'h039: dout <=  'sd1390; // 57
        'h03a: dout <=  'sd768; // 58
        'h03b: dout <=  'sd1514; // 59
        'h03c: dout <=  'sd1805; // 60
        'h03d: dout <=  'sd1536; // 61
        'h03e: dout <= -'sd1066; // 62
        'h03f: dout <= -'sd927; // 63
        'h040: dout <= -'sd1067; // 64
        'h041: dout <=  'sd2095; // 65
        'h042: dout <=  'sd1631; // 66
        'h043: dout <=  'sd2066; // 67
        'h044: dout <= -'sd1291; // 68
        'h045: dout <=  'sd1105; // 69
        'h046: dout <= -'sd2073; // 70
        'h047: dout <=  'sd402; // 71
        'h048: dout <=  'sd786; // 72
        'h049: dout <=  'sd755; // 73
        'h04a: dout <= -'sd1064; // 74
        'h04b: dout <= -'sd1272; // 75
        'h04c: dout <= -'sd766; // 76
        'h04d: dout <= -'sd2102; // 77
        'h04e: dout <=  'sd344; // 78
        'h04f: dout <= -'sd752; // 79
        'h050: dout <= -'sd1571; // 80
        'h051: dout <= -'sd1544; // 81
        'h052: dout <=  'sd919; // 82
        'h053: dout <= -'sd1323; // 83
        'h054: dout <=  'sd652; // 84
        'h055: dout <=  'sd1937; // 85
        'h056: dout <= -'sd2270; // 86
        'h057: dout <= -'sd1842; // 87
        'h058: dout <=  'sd1208; // 88
        'h059: dout <=  'sd686; // 89
        'h05a: dout <=  'sd227; // 90
        'h05b: dout <= -'sd1185; // 91
        'h05c: dout <= -'sd1492; // 92
        'h05d: dout <=  'sd1791; // 93
        'h05e: dout <=  'sd2293; // 94
        'h05f: dout <=  'sd653; // 95
        'h060: dout <= -'sd1102; // 96
        'h061: dout <=  'sd1753; // 97
        'h062: dout <=  'sd1353; // 98
        'h063: dout <= -'sd508; // 99
        'h064: dout <=  'sd1586; // 100
        'h065: dout <=  'sd1819; // 101
        'h066: dout <=  'sd81; // 102
        'h067: dout <=  'sd835; // 103
        'h068: dout <=  'sd1197; // 104
        'h069: dout <=  'sd908; // 105
        'h06a: dout <=  'sd1905; // 106
        'h06b: dout <= -'sd2108; // 107
        'h06c: dout <=  'sd1319; // 108
        'h06d: dout <= -'sd1093; // 109
        'h06e: dout <=  'sd947; // 110
        'h06f: dout <= -'sd1370; // 111
        'h070: dout <= -'sd1992; // 112
        'h071: dout <= -'sd90; // 113
        'h072: dout <= -'sd1463; // 114
        'h073: dout <= -'sd1746; // 115
        'h074: dout <= -'sd315; // 116
        'h075: dout <= -'sd1825; // 117
        'h076: dout <=  'sd116; // 118
        'h077: dout <=  'sd267; // 119
        'h078: dout <= -'sd1141; // 120
        'h079: dout <=  'sd529; // 121
        'h07a: dout <=  'sd955; // 122
        'h07b: dout <=  'sd1708; // 123
        'h07c: dout <=  'sd2045; // 124
        'h07d: dout <= -'sd2078; // 125
        'h07e: dout <= -'sd343; // 126
        'h07f: dout <= -'sd325; // 127
        'h080: dout <=  'sd673; // 128
        'h081: dout <= -'sd2098; // 129
        'h082: dout <= -'sd212; // 130
        'h083: dout <=  'sd1024; // 131
        'h084: dout <=  'sd392; // 132
        'h085: dout <=  'sd693; // 133
        'h086: dout <=  'sd599; // 134
        'h087: dout <=  'sd2193; // 135
        'h088: dout <=  'sd1112; // 136
        'h089: dout <= -'sd662; // 137
        'h08a: dout <=  'sd717; // 138
        'h08b: dout <= -'sd2175; // 139
        'h08c: dout <=  'sd1455; // 140
        'h08d: dout <=  'sd686; // 141
        'h08e: dout <=  'sd2245; // 142
        'h08f: dout <= -'sd942; // 143
        'h090: dout <=  'sd1106; // 144
        'h091: dout <=  'sd894; // 145
        'h092: dout <=  'sd1732; // 146
        'h093: dout <= -'sd1371; // 147
        'h094: dout <= -'sd1136; // 148
        'h095: dout <= -'sd1568; // 149
        'h096: dout <= -'sd960; // 150
        'h097: dout <=  'sd1319; // 151
        'h098: dout <=  'sd1215; // 152
        'h099: dout <= -'sd113; // 153
        'h09a: dout <=  'sd52; // 154
        'h09b: dout <=  'sd909; // 155
        'h09c: dout <=  'sd1098; // 156
        'h09d: dout <=  'sd167; // 157
        'h09e: dout <=  'sd1532; // 158
        'h09f: dout <= -'sd1739; // 159
        'h0a0: dout <=  'sd890; // 160
        'h0a1: dout <=  'sd960; // 161
        'h0a2: dout <= -'sd353; // 162
        'h0a3: dout <= -'sd1626; // 163
        'h0a4: dout <= -'sd415; // 164
        'h0a5: dout <=  'sd1573; // 165
        'h0a6: dout <=  'sd256; // 166
        'h0a7: dout <= -'sd512; // 167
        'h0a8: dout <=  'sd129; // 168
        'h0a9: dout <= -'sd1283; // 169
        'h0aa: dout <= -'sd1388; // 170
        'h0ab: dout <= -'sd1309; // 171
        'h0ac: dout <=  'sd2056; // 172
        'h0ad: dout <=  'sd1099; // 173
        'h0ae: dout <= -'sd2217; // 174
        'h0af: dout <= -'sd1536; // 175
        'h0b0: dout <=  'sd1585; // 176
        'h0b1: dout <= -'sd1217; // 177
        'h0b2: dout <= -'sd1591; // 178
        'h0b3: dout <=  'sd1441; // 179
        'h0b4: dout <=  'sd1287; // 180
        'h0b5: dout <= -'sd1589; // 181
        'h0b6: dout <=  'sd1498; // 182
        'h0b7: dout <= -'sd27; // 183
        'h0b8: dout <=  'sd692; // 184
        'h0b9: dout <=  'sd1372; // 185
        'h0ba: dout <= -'sd1497; // 186
        'h0bb: dout <=  'sd2190; // 187
        'h0bc: dout <= -'sd249; // 188
        'h0bd: dout <= -'sd800; // 189
        'h0be: dout <= -'sd1935; // 190
        'h0bf: dout <=  'sd1004; // 191
        'h0c0: dout <=  'sd2056; // 192
        'h0c1: dout <= -'sd2067; // 193
        'h0c2: dout <= -'sd1386; // 194
        'h0c3: dout <=  'sd1215; // 195
        'h0c4: dout <= -'sd1276; // 196
        'h0c5: dout <=  'sd510; // 197
        'h0c6: dout <=  'sd1002; // 198
        'h0c7: dout <= -'sd2228; // 199
        'h0c8: dout <= -'sd1024; // 200
        'h0c9: dout <= -'sd944; // 201
        'h0ca: dout <= -'sd2052; // 202
        'h0cb: dout <= -'sd1313; // 203
        'h0cc: dout <=  'sd2001; // 204
        'h0cd: dout <=  'sd1473; // 205
        'h0ce: dout <=  'sd1836; // 206
        'h0cf: dout <= -'sd1256; // 207
        'h0d0: dout <= -'sd584; // 208
        'h0d1: dout <=  'sd1061; // 209
        'h0d2: dout <=  'sd1222; // 210
        'h0d3: dout <= -'sd1771; // 211
        'h0d4: dout <=  'sd1662; // 212
        'h0d5: dout <= -'sd1685; // 213
        'h0d6: dout <= -'sd1090; // 214
        'h0d7: dout <=  'sd572; // 215
        'h0d8: dout <=  'sd43; // 216
        'h0d9: dout <= -'sd811; // 217
        'h0da: dout <= -'sd2036; // 218
        'h0db: dout <= -'sd278; // 219
        'h0dc: dout <=  'sd1315; // 220
        'h0dd: dout <= -'sd2015; // 221
        'h0de: dout <= -'sd911; // 222
        'h0df: dout <= -'sd248; // 223
        'h0e0: dout <=  'sd551; // 224
        'h0e1: dout <=  'sd837; // 225
        'h0e2: dout <=  'sd1307; // 226
        'h0e3: dout <= -'sd1485; // 227
        'h0e4: dout <=  'sd1345; // 228
        'h0e5: dout <= -'sd1623; // 229
        'h0e6: dout <= -'sd461; // 230
        'h0e7: dout <= -'sd1458; // 231
        'h0e8: dout <= -'sd1811; // 232
        'h0e9: dout <= -'sd1562; // 233
        'h0ea: dout <= -'sd2093; // 234
        'h0eb: dout <= -'sd1740; // 235
        'h0ec: dout <= -'sd751; // 236
        'h0ed: dout <= -'sd852; // 237
        'h0ee: dout <= -'sd19; // 238
        'h0ef: dout <= -'sd650; // 239
        'h0f0: dout <= -'sd786; // 240
        'h0f1: dout <= -'sd128; // 241
        'h0f2: dout <=  'sd1745; // 242
        'h0f3: dout <= -'sd134; // 243
        'h0f4: dout <=  'sd601; // 244
        'h0f5: dout <=  'sd2207; // 245
        'h0f6: dout <= -'sd261; // 246
        'h0f7: dout <= -'sd344; // 247
        'h0f8: dout <=  'sd872; // 248
        'h0f9: dout <= -'sd77; // 249
        'h0fa: dout <= -'sd1609; // 250
        'h0fb: dout <=  'sd905; // 251
        'h0fc: dout <= -'sd605; // 252
        'h0fd: dout <=  'sd1397; // 253
        'h0fe: dout <=  'sd1409; // 254
        'h0ff: dout <= -'sd1804; // 255
        'h100: dout <= -'sd737; // 256
        'h101: dout <=  'sd535; // 257
        'h102: dout <=  'sd249; // 258
        'h103: dout <=  'sd550; // 259
        'h104: dout <= -'sd1458; // 260
        'h105: dout <=  'sd59; // 261
        'h106: dout <=  'sd56; // 262
        'h107: dout <= -'sd1518; // 263
        'h108: dout <= -'sd1469; // 264
        'h109: dout <= -'sd2136; // 265
        'h10a: dout <=  'sd283; // 266
        'h10b: dout <=  'sd1606; // 267
        'h10c: dout <= -'sd692; // 268
        'h10d: dout <=  'sd455; // 269
        'h10e: dout <=  'sd1547; // 270
        'h10f: dout <= -'sd2125; // 271
        'h110: dout <= -'sd441; // 272
        'h111: dout <= -'sd319; // 273
        'h112: dout <=  'sd711; // 274
        'h113: dout <=  'sd34; // 275
        'h114: dout <= -'sd1223; // 276
        'h115: dout <= -'sd819; // 277
        'h116: dout <= -'sd956; // 278
        'h117: dout <=  'sd616; // 279
        'h118: dout <=  'sd810; // 280
        'h119: dout <= -'sd1308; // 281
        'h11a: dout <=  'sd1030; // 282
        'h11b: dout <=  'sd651; // 283
        'h11c: dout <=  'sd507; // 284
        'h11d: dout <= -'sd1910; // 285
        'h11e: dout <= -'sd379; // 286
        'h11f: dout <=  'sd2283; // 287
        'h120: dout <= -'sd1125; // 288
        'h121: dout <=  'sd274; // 289
        'h122: dout <= -'sd814; // 290
        'h123: dout <= -'sd1423; // 291
        'h124: dout <=  'sd927; // 292
        'h125: dout <=  'sd1083; // 293
        'h126: dout <=  'sd40; // 294
        'h127: dout <= -'sd122; // 295
        'h128: dout <=  'sd1817; // 296
        'h129: dout <= -'sd23; // 297
        'h12a: dout <=  'sd1553; // 298
        'h12b: dout <=  'sd780; // 299
        'h12c: dout <= -'sd1998; // 300
        'h12d: dout <= -'sd1612; // 301
        'h12e: dout <= -'sd34; // 302
        'h12f: dout <= -'sd511; // 303
        'h130: dout <=  'sd2118; // 304
        'h131: dout <= -'sd1750; // 305
        'h132: dout <= -'sd844; // 306
        'h133: dout <= -'sd1140; // 307
        'h134: dout <= -'sd155; // 308
        'h135: dout <=  'sd649; // 309
        'h136: dout <=  'sd1635; // 310
        'h137: dout <=  'sd2013; // 311
        'h138: dout <= -'sd96; // 312
        'h139: dout <=  'sd350; // 313
        'h13a: dout <=  'sd1743; // 314
        'h13b: dout <=  'sd298; // 315
        'h13c: dout <= -'sd126; // 316
        'h13d: dout <=  'sd1936; // 317
        'h13e: dout <= -'sd973; // 318
        'h13f: dout <=  'sd583; // 319
        'h140: dout <=  'sd2136; // 320
        'h141: dout <=  'sd2194; // 321
        'h142: dout <= -'sd1724; // 322
        'h143: dout <= -'sd2083; // 323
        'h144: dout <=  'sd875; // 324
        'h145: dout <=  'sd1860; // 325
        'h146: dout <= -'sd1697; // 326
        'h147: dout <=  'sd1473; // 327
        'h148: dout <=  'sd107; // 328
        'h149: dout <= -'sd2148; // 329
        'h14a: dout <= -'sd2273; // 330
        'h14b: dout <=  'sd2204; // 331
        'h14c: dout <=  'sd335; // 332
        'h14d: dout <=  'sd707; // 333
        'h14e: dout <= -'sd42; // 334
        'h14f: dout <= -'sd561; // 335
        'h150: dout <=  'sd2244; // 336
        'h151: dout <=  'sd1466; // 337
        'h152: dout <=  'sd1573; // 338
        'h153: dout <= -'sd1767; // 339
        'h154: dout <= -'sd2150; // 340
        'h155: dout <=  'sd1416; // 341
        'h156: dout <= -'sd2032; // 342
        'h157: dout <= -'sd1119; // 343
        'h158: dout <=  'sd1824; // 344
        'h159: dout <= -'sd353; // 345
        'h15a: dout <=  'sd1990; // 346
        'h15b: dout <= -'sd48; // 347
        'h15c: dout <=  'sd743; // 348
        'h15d: dout <=  'sd1089; // 349
        'h15e: dout <=  'sd1982; // 350
        'h15f: dout <=  'sd1830; // 351
        'h160: dout <= -'sd1533; // 352
        'h161: dout <=  'sd2057; // 353
        'h162: dout <=  'sd1039; // 354
        'h163: dout <=  'sd367; // 355
        'h164: dout <= -'sd2229; // 356
        'h165: dout <=  'sd651; // 357
        'h166: dout <= -'sd1493; // 358
        'h167: dout <=  'sd1459; // 359
        'h168: dout <=  'sd691; // 360
        'h169: dout <= -'sd861; // 361
        'h16a: dout <=  'sd2202; // 362
        'h16b: dout <= -'sd619; // 363
        'h16c: dout <=  'sd804; // 364
        'h16d: dout <=  'sd1927; // 365
        'h16e: dout <= -'sd2203; // 366
        'h16f: dout <=  'sd2139; // 367
        'h170: dout <= -'sd1426; // 368
        'h171: dout <= -'sd2053; // 369
        'h172: dout <= -'sd2216; // 370
        'h173: dout <=  'sd1074; // 371
        'h174: dout <=  'sd1007; // 372
        'h175: dout <=  'sd1580; // 373
        'h176: dout <=  'sd2034; // 374
        'h177: dout <= -'sd176; // 375
        'h178: dout <= -'sd1812; // 376
        'h179: dout <=  'sd2151; // 377
        'h17a: dout <=  'sd1774; // 378
        'h17b: dout <= -'sd2072; // 379
        'h17c: dout <=  'sd1532; // 380
        'h17d: dout <=  'sd2271; // 381
        'h17e: dout <= -'sd995; // 382
        'h17f: dout <=  'sd28; // 383
        'h180: dout <=  'sd1883; // 384
        'h181: dout <=  'sd223; // 385
        'h182: dout <= -'sd190; // 386
        'h183: dout <=  'sd714; // 387
        'h184: dout <=  'sd2052; // 388
        'h185: dout <= -'sd831; // 389
        'h186: dout <=  'sd616; // 390
        'h187: dout <=  'sd1789; // 391
        'h188: dout <=  'sd1216; // 392
        'h189: dout <=  'sd1728; // 393
        'h18a: dout <=  'sd1923; // 394
        'h18b: dout <=  'sd447; // 395
        'h18c: dout <= -'sd446; // 396
        'h18d: dout <=  'sd2241; // 397
        'h18e: dout <= -'sd565; // 398
        'h18f: dout <= -'sd1456; // 399
        'h190: dout <= -'sd1798; // 400
        'h191: dout <= -'sd846; // 401
        'h192: dout <=  'sd1099; // 402
        'h193: dout <=  'sd47; // 403
        'h194: dout <=  'sd1137; // 404
        'h195: dout <= -'sd482; // 405
        'h196: dout <=  'sd37; // 406
        'h197: dout <=  'sd1252; // 407
        'h198: dout <=  'sd1671; // 408
        'h199: dout <=  'sd1317; // 409
        'h19a: dout <=  'sd675; // 410
        'h19b: dout <=  'sd0; // 411
        'h19c: dout <= -'sd554; // 412
        'h19d: dout <= -'sd983; // 413
        'h19e: dout <= -'sd839; // 414
        'h19f: dout <= -'sd2059; // 415
        'h1a0: dout <= -'sd199; // 416
        'h1a1: dout <=  'sd1031; // 417
        'h1a2: dout <=  'sd1026; // 418
        'h1a3: dout <= -'sd308; // 419
        'h1a4: dout <= -'sd186; // 420
        'h1a5: dout <= -'sd1271; // 421
        'h1a6: dout <= -'sd378; // 422
        'h1a7: dout <=  'sd2128; // 423
        'h1a8: dout <= -'sd599; // 424
        'h1a9: dout <=  'sd1317; // 425
        'h1aa: dout <=  'sd719; // 426
        'h1ab: dout <= -'sd224; // 427
        'h1ac: dout <= -'sd1763; // 428
        'h1ad: dout <= -'sd1378; // 429
        'h1ae: dout <= -'sd1446; // 430
        'h1af: dout <= -'sd1748; // 431
        'h1b0: dout <= -'sd1299; // 432
        'h1b1: dout <= -'sd265; // 433
        'h1b2: dout <=  'sd2196; // 434
        'h1b3: dout <= -'sd1851; // 435
        'h1b4: dout <= -'sd2258; // 436
        'h1b5: dout <=  'sd1240; // 437
        'h1b6: dout <= -'sd221; // 438
        'h1b7: dout <= -'sd1463; // 439
        'h1b8: dout <=  'sd484; // 440
        'h1b9: dout <=  'sd742; // 441
        'h1ba: dout <= -'sd517; // 442
        'h1bb: dout <= -'sd2198; // 443
        'h1bc: dout <= -'sd402; // 444
        'h1bd: dout <= -'sd1236; // 445
        'h1be: dout <= -'sd1327; // 446
        'h1bf: dout <= -'sd1849; // 447
        'h1c0: dout <= -'sd1613; // 448
        'h1c1: dout <= -'sd1368; // 449
        'h1c2: dout <= -'sd1191; // 450
        'h1c3: dout <=  'sd402; // 451
        'h1c4: dout <=  'sd332; // 452
        'h1c5: dout <= -'sd838; // 453
        'h1c6: dout <= -'sd1948; // 454
        'h1c7: dout <= -'sd824; // 455
        'h1c8: dout <= -'sd1887; // 456
        'h1c9: dout <=  'sd1469; // 457
        'h1ca: dout <= -'sd1950; // 458
        'h1cb: dout <=  'sd1153; // 459
        'h1cc: dout <=  'sd1218; // 460
        'h1cd: dout <= -'sd1362; // 461
        'h1ce: dout <=  'sd23; // 462
        'h1cf: dout <= -'sd1370; // 463
        'h1d0: dout <=  'sd142; // 464
        'h1d1: dout <=  'sd460; // 465
        'h1d2: dout <= -'sd1140; // 466
        'h1d3: dout <= -'sd1491; // 467
        'h1d4: dout <= -'sd490; // 468
        'h1d5: dout <=  'sd2221; // 469
        'h1d6: dout <= -'sd1438; // 470
        'h1d7: dout <=  'sd1191; // 471
        'h1d8: dout <= -'sd2292; // 472
        'h1d9: dout <=  'sd1148; // 473
        'h1da: dout <=  'sd378; // 474
        'h1db: dout <= -'sd2016; // 475
        'h1dc: dout <=  'sd1951; // 476
        'h1dd: dout <=  'sd3; // 477
        'h1de: dout <=  'sd1278; // 478
        'h1df: dout <= -'sd20; // 479
        'h1e0: dout <= -'sd1843; // 480
        'h1e1: dout <=  'sd2234; // 481
        'h1e2: dout <=  'sd276; // 482
        'h1e3: dout <=  'sd1739; // 483
        'h1e4: dout <= -'sd1895; // 484
        'h1e5: dout <=  'sd29; // 485
        'h1e6: dout <=  'sd2241; // 486
        'h1e7: dout <=  'sd466; // 487
        'h1e8: dout <=  'sd308; // 488
        'h1e9: dout <=  'sd571; // 489
        'h1ea: dout <=  'sd612; // 490
        'h1eb: dout <=  'sd1495; // 491
        'h1ec: dout <= -'sd706; // 492
        'h1ed: dout <= -'sd2026; // 493
        'h1ee: dout <= -'sd1213; // 494
        'h1ef: dout <=  'sd604; // 495
        'h1f0: dout <= -'sd91; // 496
        'h1f1: dout <= -'sd2293; // 497
        'h1f2: dout <= -'sd390; // 498
        'h1f3: dout <=  'sd374; // 499
        'h1f4: dout <= -'sd691; // 500
        'h1f5: dout <=  'sd2146; // 501
        'h1f6: dout <= -'sd1342; // 502
        'h1f7: dout <= -'sd870; // 503
        'h1f8: dout <= -'sd215; // 504
        'h1f9: dout <= -'sd2042; // 505
        'h1fa: dout <= -'sd450; // 506
        'h1fb: dout <= -'sd2260; // 507
        'h1fc: dout <=  'sd629; // 508
        'h1fd: dout <= -'sd1787; // 509
        'h1fe: dout <= -'sd2066; // 510
        'h1ff: dout <=  'sd1603; // 511
        'h200: dout <=  'sd1050; // 512
        'h201: dout <= -'sd1379; // 513
        'h202: dout <=  'sd1393; // 514
        'h203: dout <=  'sd390; // 515
        'h204: dout <=  'sd1082; // 516
        'h205: dout <=  'sd488; // 517
        'h206: dout <=  'sd892; // 518
        'h207: dout <= -'sd163; // 519
        'h208: dout <=  'sd310; // 520
        'h209: dout <=  'sd1382; // 521
        'h20a: dout <=  'sd104; // 522
        'h20b: dout <=  'sd696; // 523
        'h20c: dout <=  'sd2041; // 524
        'h20d: dout <= -'sd157; // 525
        'h20e: dout <=  'sd567; // 526
        'h20f: dout <=  'sd189; // 527
        'h210: dout <=  'sd268; // 528
        'h211: dout <= -'sd1148; // 529
        'h212: dout <=  'sd310; // 530
        'h213: dout <= -'sd760; // 531
        'h214: dout <=  'sd2051; // 532
        'h215: dout <=  'sd464; // 533
        'h216: dout <=  'sd977; // 534
        'h217: dout <= -'sd1294; // 535
        'h218: dout <=  'sd1373; // 536
        'h219: dout <= -'sd1137; // 537
        'h21a: dout <= -'sd1178; // 538
        'h21b: dout <= -'sd2177; // 539
        'h21c: dout <=  'sd2228; // 540
        'h21d: dout <=  'sd1777; // 541
        'h21e: dout <= -'sd1468; // 542
        'h21f: dout <=  'sd1224; // 543
        'h220: dout <=  'sd1161; // 544
        'h221: dout <= -'sd1090; // 545
        'h222: dout <= -'sd1069; // 546
        'h223: dout <=  'sd238; // 547
        'h224: dout <= -'sd976; // 548
        'h225: dout <=  'sd1655; // 549
        'h226: dout <=  'sd205; // 550
        'h227: dout <=  'sd1989; // 551
        'h228: dout <= -'sd1850; // 552
        'h229: dout <= -'sd817; // 553
        'h22a: dout <=  'sd475; // 554
        'h22b: dout <=  'sd1322; // 555
        'h22c: dout <=  'sd596; // 556
        'h22d: dout <=  'sd1970; // 557
        'h22e: dout <= -'sd424; // 558
        'h22f: dout <=  'sd409; // 559
        'h230: dout <= -'sd647; // 560
        'h231: dout <=  'sd941; // 561
        'h232: dout <= -'sd2189; // 562
        'h233: dout <=  'sd683; // 563
        'h234: dout <=  'sd1880; // 564
        'h235: dout <= -'sd90; // 565
        'h236: dout <=  'sd1207; // 566
        'h237: dout <= -'sd1018; // 567
        'h238: dout <= -'sd2224; // 568
        'h239: dout <=  'sd511; // 569
        'h23a: dout <= -'sd58; // 570
        'h23b: dout <= -'sd877; // 571
        'h23c: dout <= -'sd2037; // 572
        'h23d: dout <= -'sd1486; // 573
        'h23e: dout <=  'sd1739; // 574
        'h23f: dout <=  'sd159; // 575
        'h240: dout <= -'sd971; // 576
        'h241: dout <=  'sd1848; // 577
        'h242: dout <=  'sd79; // 578
        'h243: dout <= -'sd1141; // 579
        'h244: dout <= -'sd1296; // 580
        'h245: dout <= -'sd29; // 581
        'h246: dout <= -'sd712; // 582
        'h247: dout <= -'sd145; // 583
        'h248: dout <=  'sd85; // 584
        'h249: dout <= -'sd945; // 585
        'h24a: dout <=  'sd398; // 586
        'h24b: dout <=  'sd662; // 587
        'h24c: dout <= -'sd743; // 588
        'h24d: dout <=  'sd660; // 589
        'h24e: dout <= -'sd219; // 590
        'h24f: dout <= -'sd882; // 591
        'h250: dout <= -'sd1584; // 592
        'h251: dout <=  'sd1132; // 593
        'h252: dout <= -'sd561; // 594
        'h253: dout <= -'sd534; // 595
        'h254: dout <= -'sd747; // 596
        'h255: dout <= -'sd1263; // 597
        'h256: dout <= -'sd367; // 598
        'h257: dout <=  'sd1630; // 599
        'h258: dout <=  'sd390; // 600
        'h259: dout <=  'sd1276; // 601
        'h25a: dout <=  'sd1715; // 602
        'h25b: dout <= -'sd1970; // 603
        'h25c: dout <=  'sd80; // 604
        'h25d: dout <= -'sd1913; // 605
        'h25e: dout <=  'sd19; // 606
        'h25f: dout <=  'sd2144; // 607
        'h260: dout <= -'sd1810; // 608
        'h261: dout <= -'sd1241; // 609
        'h262: dout <= -'sd2245; // 610
        'h263: dout <=  'sd648; // 611
        'h264: dout <=  'sd474; // 612
        'h265: dout <=  'sd1690; // 613
        'h266: dout <= -'sd682; // 614
        'h267: dout <= -'sd2057; // 615
        'h268: dout <= -'sd1211; // 616
        'h269: dout <=  'sd533; // 617
        'h26a: dout <=  'sd1971; // 618
        'h26b: dout <=  'sd895; // 619
        'h26c: dout <= -'sd1269; // 620
        'h26d: dout <= -'sd614; // 621
        'h26e: dout <=  'sd2038; // 622
        'h26f: dout <= -'sd1752; // 623
        'h270: dout <= -'sd282; // 624
        'h271: dout <= -'sd884; // 625
        'h272: dout <= -'sd1689; // 626
        'h273: dout <= -'sd1292; // 627
        'h274: dout <= -'sd801; // 628
        'h275: dout <=  'sd1529; // 629
        'h276: dout <= -'sd486; // 630
        'h277: dout <= -'sd1990; // 631
        'h278: dout <=  'sd1041; // 632
        'h279: dout <=  'sd195; // 633
        'h27a: dout <=  'sd885; // 634
        'h27b: dout <=  'sd105; // 635
        'h27c: dout <= -'sd1136; // 636
        'h27d: dout <=  'sd187; // 637
        'h27e: dout <=  'sd395; // 638
        'h27f: dout <= -'sd2; // 639
        'h280: dout <= -'sd868; // 640
        'h281: dout <= -'sd1454; // 641
        'h282: dout <=  'sd50; // 642
        'h283: dout <= -'sd831; // 643
        'h284: dout <=  'sd1728; // 644
        'h285: dout <= -'sd1416; // 645
        'h286: dout <= -'sd1220; // 646
        'h287: dout <= -'sd2270; // 647
        'h288: dout <=  'sd1533; // 648
        'h289: dout <=  'sd1256; // 649
        'h28a: dout <= -'sd3; // 650
        'h28b: dout <=  'sd64; // 651
        'h28c: dout <= -'sd472; // 652
        'h28d: dout <=  'sd622; // 653
        'h28e: dout <= -'sd232; // 654
        'h28f: dout <= -'sd64; // 655
        'h290: dout <= -'sd2174; // 656
        'h291: dout <= -'sd820; // 657
        'h292: dout <= -'sd184; // 658
        'h293: dout <= -'sd2285; // 659
        'h294: dout <=  'sd717; // 660
        'h295: dout <=  'sd353; // 661
        'h296: dout <=  'sd2103; // 662
        'h297: dout <=  'sd228; // 663
        'h298: dout <=  'sd472; // 664
        'h299: dout <= -'sd698; // 665
        'h29a: dout <= -'sd949; // 666
        'h29b: dout <=  'sd361; // 667
        'h29c: dout <=  'sd1096; // 668
        'h29d: dout <=  'sd1160; // 669
        'h29e: dout <=  'sd2111; // 670
        'h29f: dout <=  'sd2; // 671
        'h2a0: dout <=  'sd1620; // 672
        'h2a1: dout <=  'sd1041; // 673
        'h2a2: dout <=  'sd1313; // 674
        'h2a3: dout <= -'sd206; // 675
        'h2a4: dout <= -'sd657; // 676
        'h2a5: dout <= -'sd2144; // 677
        'h2a6: dout <= -'sd2171; // 678
        'h2a7: dout <= -'sd1296; // 679
        'h2a8: dout <= -'sd1489; // 680
        'h2a9: dout <= -'sd1155; // 681
        'h2aa: dout <= -'sd649; // 682
        'h2ab: dout <=  'sd1308; // 683
        'h2ac: dout <= -'sd2089; // 684
        'h2ad: dout <=  'sd475; // 685
        'h2ae: dout <=  'sd237; // 686
        'h2af: dout <= -'sd1124; // 687
        'h2b0: dout <= -'sd874; // 688
        'h2b1: dout <=  'sd47; // 689
        'h2b2: dout <= -'sd501; // 690
        'h2b3: dout <= -'sd2010; // 691
        'h2b4: dout <= -'sd62; // 692
        'h2b5: dout <= -'sd1462; // 693
        'h2b6: dout <=  'sd205; // 694
        'h2b7: dout <= -'sd105; // 695
        'h2b8: dout <= -'sd831; // 696
        'h2b9: dout <=  'sd2152; // 697
        'h2ba: dout <= -'sd1827; // 698
        'h2bb: dout <= -'sd1070; // 699
        'h2bc: dout <=  'sd1780; // 700
        'h2bd: dout <=  'sd292; // 701
        'h2be: dout <=  'sd1623; // 702
        'h2bf: dout <= -'sd2060; // 703
        'h2c0: dout <= -'sd716; // 704
        'h2c1: dout <=  'sd204; // 705
        'h2c2: dout <=  'sd718; // 706
        'h2c3: dout <=  'sd832; // 707
        'h2c4: dout <=  'sd1724; // 708
        'h2c5: dout <=  'sd99; // 709
        'h2c6: dout <=  'sd1813; // 710
        'h2c7: dout <= -'sd924; // 711
        'h2c8: dout <= -'sd1215; // 712
        'h2c9: dout <=  'sd2278; // 713
        'h2ca: dout <= -'sd85; // 714
        'h2cb: dout <= -'sd791; // 715
        'h2cc: dout <=  'sd2280; // 716
        'h2cd: dout <=  'sd1032; // 717
        'h2ce: dout <=  'sd1680; // 718
        'h2cf: dout <= -'sd140; // 719
        'h2d0: dout <=  'sd550; // 720
        'h2d1: dout <= -'sd1608; // 721
        'h2d2: dout <= -'sd1488; // 722
        'h2d3: dout <=  'sd1005; // 723
        'h2d4: dout <= -'sd272; // 724
        'h2d5: dout <=  'sd681; // 725
        'h2d6: dout <= -'sd202; // 726
        'h2d7: dout <= -'sd1667; // 727
        'h2d8: dout <=  'sd1860; // 728
        'h2d9: dout <=  'sd549; // 729
        'h2da: dout <=  'sd1268; // 730
        'h2db: dout <=  'sd1358; // 731
        'h2dc: dout <= -'sd1066; // 732
        'h2dd: dout <=  'sd132; // 733
        'h2de: dout <= -'sd2038; // 734
        'h2df: dout <= -'sd810; // 735
        'h2e0: dout <=  'sd2229; // 736
        'h2e1: dout <= -'sd1555; // 737
        'h2e2: dout <= -'sd906; // 738
        'h2e3: dout <=  'sd59; // 739
        'h2e4: dout <=  'sd1439; // 740
        'h2e5: dout <= -'sd1673; // 741
        'h2e6: dout <= -'sd29; // 742
        'h2e7: dout <= -'sd1060; // 743
        'h2e8: dout <=  'sd1968; // 744
        'h2e9: dout <= -'sd1516; // 745
        'h2ea: dout <=  'sd501; // 746
        'h2eb: dout <= -'sd896; // 747
        'h2ec: dout <=  'sd1882; // 748
        'h2ed: dout <= -'sd292; // 749
        'h2ee: dout <=  'sd1798; // 750
        'h2ef: dout <= -'sd1682; // 751
        'h2f0: dout <= -'sd106; // 752
        'h2f1: dout <=  'sd1069; // 753
        'h2f2: dout <=  'sd1227; // 754
        'h2f3: dout <=  'sd236; // 755
        'h2f4: dout <=  'sd1347; // 756
        'h2f5: dout <=  'sd2120; // 757
        'h2f6: dout <= -'sd151; // 758
        'h2f7: dout <= -'sd994; // 759
        'h2f8: dout <=  'sd2212; // 760
        'h2f9: dout <=  'sd869; // 761
        'h2fa: dout <=  'sd1492; // 762
        'h2fb: dout <=  'sd1827; // 763
        'h2fc: dout <= -'sd1248; // 764
        'h2fd: dout <=  'sd1372; // 765
        'h2fe: dout <=  'sd555; // 766
        'h2ff: dout <= -'sd169; // 767
        'h300: dout <= -'sd2108; // 768
        'h301: dout <=  'sd969; // 769
        'h302: dout <= -'sd34; // 770
        'h303: dout <= -'sd1453; // 771
        'h304: dout <= -'sd425; // 772
        'h305: dout <= -'sd596; // 773
        'h306: dout <=  'sd1287; // 774
        'h307: dout <= -'sd35; // 775
        'h308: dout <= -'sd993; // 776
        'h309: dout <= -'sd1080; // 777
        'h30a: dout <= -'sd71; // 778
        'h30b: dout <= -'sd2171; // 779
        'h30c: dout <=  'sd1205; // 780
        'h30d: dout <=  'sd1994; // 781
        'h30e: dout <= -'sd1411; // 782
        'h30f: dout <= -'sd1730; // 783
        'h310: dout <= -'sd2265; // 784
        'h311: dout <=  'sd56; // 785
        'h312: dout <= -'sd2165; // 786
        'h313: dout <=  'sd1644; // 787
        'h314: dout <= -'sd1965; // 788
        'h315: dout <=  'sd1527; // 789
        'h316: dout <=  'sd1431; // 790
        'h317: dout <= -'sd1087; // 791
        'h318: dout <= -'sd998; // 792
        'h319: dout <=  'sd2090; // 793
        'h31a: dout <= -'sd1960; // 794
        'h31b: dout <=  'sd691; // 795
        'h31c: dout <= -'sd447; // 796
        'h31d: dout <= -'sd1854; // 797
        'h31e: dout <=  'sd1046; // 798
        'h31f: dout <=  'sd35; // 799
        'h320: dout <= -'sd613; // 800
        'h321: dout <= -'sd1826; // 801
        'h322: dout <=  'sd1831; // 802
        'h323: dout <=  'sd1098; // 803
        'h324: dout <= -'sd1518; // 804
        'h325: dout <=  'sd562; // 805
        'h326: dout <= -'sd1317; // 806
        'h327: dout <= -'sd682; // 807
        'h328: dout <=  'sd818; // 808
        'h329: dout <= -'sd2158; // 809
        'h32a: dout <= -'sd404; // 810
        'h32b: dout <= -'sd1418; // 811
        'h32c: dout <=  'sd1838; // 812
        'h32d: dout <=  'sd377; // 813
        'h32e: dout <= -'sd778; // 814
        'h32f: dout <= -'sd126; // 815
        'h330: dout <=  'sd1615; // 816
        'h331: dout <= -'sd1361; // 817
        'h332: dout <= -'sd1634; // 818
        'h333: dout <= -'sd2068; // 819
        'h334: dout <=  'sd1975; // 820
        'h335: dout <=  'sd950; // 821
        'h336: dout <=  'sd1858; // 822
        'h337: dout <=  'sd36; // 823
        'h338: dout <=  'sd41; // 824
        'h339: dout <=  'sd1464; // 825
        'h33a: dout <=  'sd576; // 826
        'h33b: dout <= -'sd1010; // 827
        'h33c: dout <=  'sd26; // 828
        'h33d: dout <=  'sd1447; // 829
        'h33e: dout <= -'sd220; // 830
        'h33f: dout <= -'sd1447; // 831
        'h340: dout <= -'sd1301; // 832
        'h341: dout <= -'sd467; // 833
        'h342: dout <= -'sd149; // 834
        'h343: dout <=  'sd2040; // 835
        'h344: dout <=  'sd1885; // 836
        'h345: dout <=  'sd2175; // 837
        'h346: dout <= -'sd1640; // 838
        'h347: dout <= -'sd412; // 839
        'h348: dout <=  'sd630; // 840
        'h349: dout <=  'sd1868; // 841
        'h34a: dout <=  'sd521; // 842
        'h34b: dout <= -'sd1636; // 843
        'h34c: dout <=  'sd1835; // 844
        'h34d: dout <= -'sd723; // 845
        'h34e: dout <=  'sd531; // 846
        'h34f: dout <=  'sd2063; // 847
        'h350: dout <=  'sd2250; // 848
        'h351: dout <=  'sd64; // 849
        'h352: dout <= -'sd1549; // 850
        'h353: dout <=  'sd1384; // 851
        'h354: dout <= -'sd257; // 852
        'h355: dout <=  'sd2101; // 853
        'h356: dout <=  'sd420; // 854
        'h357: dout <= -'sd2243; // 855
        'h358: dout <=  'sd1963; // 856
        'h359: dout <= -'sd1178; // 857
        'h35a: dout <= -'sd1903; // 858
        'h35b: dout <=  'sd826; // 859
        'h35c: dout <= -'sd966; // 860
        'h35d: dout <=  'sd693; // 861
        'h35e: dout <= -'sd1296; // 862
        'h35f: dout <= -'sd32; // 863
        'h360: dout <=  'sd2159; // 864
        'h361: dout <=  'sd180; // 865
        'h362: dout <=  'sd1057; // 866
        'h363: dout <=  'sd2248; // 867
        'h364: dout <=  'sd2238; // 868
        'h365: dout <=  'sd2073; // 869
        'h366: dout <= -'sd446; // 870
        'h367: dout <= -'sd452; // 871
        'h368: dout <=  'sd289; // 872
        'h369: dout <= -'sd213; // 873
        'h36a: dout <=  'sd331; // 874
        'h36b: dout <= -'sd846; // 875
        'h36c: dout <=  'sd1048; // 876
        'h36d: dout <=  'sd1048; // 877
        'h36e: dout <= -'sd769; // 878
        'h36f: dout <=  'sd498; // 879
        'h370: dout <= -'sd2039; // 880
        'h371: dout <=  'sd1669; // 881
        'h372: dout <= -'sd505; // 882
        'h373: dout <= -'sd383; // 883
        'h374: dout <= -'sd2275; // 884
        'h375: dout <=  'sd545; // 885
        'h376: dout <=  'sd2055; // 886
        'h377: dout <= -'sd1846; // 887
        'h378: dout <=  'sd1895; // 888
        'h379: dout <= -'sd1289; // 889
        'h37a: dout <=  'sd1654; // 890
        'h37b: dout <=  'sd528; // 891
        'h37c: dout <=  'sd1363; // 892
        'h37d: dout <=  'sd1635; // 893
        'h37e: dout <= -'sd1084; // 894
        'h37f: dout <=  'sd864; // 895
        'h380: dout <= -'sd1311; // 896
        'h381: dout <=  'sd1477; // 897
        'h382: dout <=  'sd178; // 898
        'h383: dout <= -'sd1986; // 899
        'h384: dout <= -'sd2059; // 900
        'h385: dout <=  'sd1614; // 901
        'h386: dout <=  'sd750; // 902
        'h387: dout <=  'sd1125; // 903
        'h388: dout <= -'sd1940; // 904
        'h389: dout <=  'sd671; // 905
        'h38a: dout <=  'sd327; // 906
        'h38b: dout <=  'sd1594; // 907
        'h38c: dout <= -'sd1670; // 908
        'h38d: dout <=  'sd1096; // 909
        'h38e: dout <= -'sd1258; // 910
        'h38f: dout <= -'sd641; // 911
        'h390: dout <= -'sd2030; // 912
        'h391: dout <=  'sd2042; // 913
        'h392: dout <=  'sd1640; // 914
        'h393: dout <=  'sd2232; // 915
        'h394: dout <=  'sd983; // 916
        'h395: dout <=  'sd2228; // 917
        'h396: dout <=  'sd32; // 918
        'h397: dout <=  'sd1033; // 919
        'h398: dout <= -'sd985; // 920
        'h399: dout <=  'sd1092; // 921
        'h39a: dout <=  'sd2041; // 922
        'h39b: dout <= -'sd2054; // 923
        'h39c: dout <=  'sd2073; // 924
        'h39d: dout <=  'sd1214; // 925
        'h39e: dout <= -'sd1301; // 926
        'h39f: dout <= -'sd2218; // 927
        'h3a0: dout <=  'sd889; // 928
        'h3a1: dout <= -'sd14; // 929
        'h3a2: dout <=  'sd1459; // 930
        'h3a3: dout <= -'sd1373; // 931
        'h3a4: dout <= -'sd1147; // 932
        'h3a5: dout <= -'sd1947; // 933
        'h3a6: dout <=  'sd212; // 934
        'h3a7: dout <= -'sd436; // 935
        'h3a8: dout <=  'sd360; // 936
        'h3a9: dout <= -'sd754; // 937
        'h3aa: dout <=  'sd2276; // 938
        'h3ab: dout <=  'sd664; // 939
        'h3ac: dout <=  'sd2156; // 940
        'h3ad: dout <=  'sd2205; // 941
        'h3ae: dout <=  'sd591; // 942
        'h3af: dout <=  'sd2152; // 943
        'h3b0: dout <=  'sd1790; // 944
        'h3b1: dout <= -'sd1265; // 945
        'h3b2: dout <= -'sd86; // 946
        'h3b3: dout <=  'sd1782; // 947
        'h3b4: dout <= -'sd198; // 948
        'h3b5: dout <= -'sd519; // 949
        'h3b6: dout <=  'sd2279; // 950
        'h3b7: dout <= -'sd1530; // 951
        'h3b8: dout <=  'sd1122; // 952
        'h3b9: dout <=  'sd495; // 953
        'h3ba: dout <= -'sd1790; // 954
        'h3bb: dout <= -'sd1013; // 955
        'h3bc: dout <= -'sd37; // 956
        'h3bd: dout <= -'sd133; // 957
        'h3be: dout <=  'sd1073; // 958
        'h3bf: dout <=  'sd944; // 959
        'h3c0: dout <=  'sd1872; // 960
        'h3c1: dout <=  'sd1568; // 961
        'h3c2: dout <= -'sd570; // 962
        'h3c3: dout <= -'sd142; // 963
        'h3c4: dout <= -'sd429; // 964
        'h3c5: dout <=  'sd873; // 965
        'h3c6: dout <= -'sd2267; // 966
        'h3c7: dout <= -'sd1430; // 967
        'h3c8: dout <=  'sd2171; // 968
        'h3c9: dout <=  'sd1339; // 969
        'h3ca: dout <=  'sd334; // 970
        'h3cb: dout <=  'sd1644; // 971
        'h3cc: dout <= -'sd1504; // 972
        'h3cd: dout <=  'sd862; // 973
        'h3ce: dout <= -'sd564; // 974
        'h3cf: dout <=  'sd846; // 975
        'h3d0: dout <= -'sd858; // 976
        'h3d1: dout <= -'sd633; // 977
        'h3d2: dout <=  'sd2003; // 978
        'h3d3: dout <= -'sd2145; // 979
        'h3d4: dout <= -'sd1495; // 980
        'h3d5: dout <= -'sd1883; // 981
        'h3d6: dout <= -'sd840; // 982
        'h3d7: dout <=  'sd1216; // 983
        'h3d8: dout <= -'sd1395; // 984
        'h3d9: dout <=  'sd211; // 985
        'h3da: dout <= -'sd1753; // 986
        'h3db: dout <= -'sd1436; // 987
        'h3dc: dout <= -'sd1008; // 988
        'h3dd: dout <=  'sd194; // 989
        'h3de: dout <= -'sd1882; // 990
        'h3df: dout <=  'sd1934; // 991
        'h3e0: dout <=  'sd533; // 992
        'h3e1: dout <=  'sd1725; // 993
        'h3e2: dout <= -'sd2255; // 994
        'h3e3: dout <=  'sd1821; // 995
        'h3e4: dout <= -'sd94; // 996
        'h3e5: dout <= -'sd612; // 997
        'h3e6: dout <= -'sd1552; // 998
        'h3e7: dout <= -'sd1495; // 999
        'h3e8: dout <= -'sd98; // 1000
        'h3e9: dout <=  'sd271; // 1001
        'h3ea: dout <= -'sd260; // 1002
        'h3eb: dout <= -'sd227; // 1003
        'h3ec: dout <= -'sd1507; // 1004
        'h3ed: dout <= -'sd1487; // 1005
        'h3ee: dout <=  'sd1894; // 1006
        'h3ef: dout <=  'sd1650; // 1007
        'h3f0: dout <=  'sd456; // 1008
        'h3f1: dout <= -'sd819; // 1009
        'h3f2: dout <= -'sd1796; // 1010
        'h3f3: dout <=  'sd491; // 1011
        'h3f4: dout <= -'sd1039; // 1012
        'h3f5: dout <= -'sd577; // 1013
        'h3f6: dout <= -'sd1271; // 1014
        'h3f7: dout <= -'sd477; // 1015
        'h3f8: dout <=  'sd110; // 1016
        'h3f9: dout <= -'sd2069; // 1017
        'h3fa: dout <=  'sd1252; // 1018
        'h3fb: dout <= -'sd2131; // 1019
        'h3fc: dout <=  'sd2285; // 1020
        'h3fd: dout <= -'sd2055; // 1021
        'h3fe: dout <= -'sd661; // 1022
        'h3ff: dout <=  'sd1412; // 1023
        'h400: dout <=  'sd2264; // 1024
        'h401: dout <=  'sd1805; // 1025
        'h402: dout <=  'sd2145; // 1026
        'h403: dout <=  'sd110; // 1027
        'h404: dout <= -'sd936; // 1028
        'h405: dout <= -'sd1648; // 1029
        'h406: dout <=  'sd229; // 1030
        'h407: dout <=  'sd1561; // 1031
        'h408: dout <= -'sd485; // 1032
        'h409: dout <= -'sd80; // 1033
        'h40a: dout <= -'sd1847; // 1034
        'h40b: dout <=  'sd179; // 1035
        'h40c: dout <= -'sd1635; // 1036
        'h40d: dout <= -'sd136; // 1037
        'h40e: dout <=  'sd1629; // 1038
        'h40f: dout <= -'sd1319; // 1039
        'h410: dout <=  'sd840; // 1040
        'h411: dout <=  'sd1399; // 1041
        'h412: dout <= -'sd1139; // 1042
        'h413: dout <=  'sd329; // 1043
        'h414: dout <= -'sd1544; // 1044
        'h415: dout <=  'sd1746; // 1045
        'h416: dout <=  'sd1620; // 1046
        'h417: dout <=  'sd239; // 1047
        'h418: dout <=  'sd2076; // 1048
        'h419: dout <= -'sd123; // 1049
        'h41a: dout <=  'sd1693; // 1050
        'h41b: dout <=  'sd503; // 1051
        'h41c: dout <=  'sd569; // 1052
        'h41d: dout <= -'sd921; // 1053
        'h41e: dout <=  'sd267; // 1054
        'h41f: dout <= -'sd1068; // 1055
        'h420: dout <=  'sd1429; // 1056
        'h421: dout <= -'sd724; // 1057
        'h422: dout <= -'sd982; // 1058
        'h423: dout <=  'sd556; // 1059
        'h424: dout <=  'sd1366; // 1060
        'h425: dout <=  'sd1486; // 1061
        'h426: dout <= -'sd617; // 1062
        'h427: dout <= -'sd2190; // 1063
        'h428: dout <=  'sd802; // 1064
        'h429: dout <= -'sd636; // 1065
        'h42a: dout <= -'sd1972; // 1066
        'h42b: dout <= -'sd2173; // 1067
        'h42c: dout <= -'sd1839; // 1068
        'h42d: dout <=  'sd2209; // 1069
        'h42e: dout <=  'sd1674; // 1070
        'h42f: dout <= -'sd1937; // 1071
        'h430: dout <= -'sd628; // 1072
        'h431: dout <= -'sd1739; // 1073
        'h432: dout <=  'sd1462; // 1074
        'h433: dout <= -'sd439; // 1075
        'h434: dout <=  'sd757; // 1076
        'h435: dout <=  'sd2280; // 1077
        'h436: dout <=  'sd1713; // 1078
        'h437: dout <= -'sd1129; // 1079
        'h438: dout <=  'sd948; // 1080
        'h439: dout <= -'sd1862; // 1081
        'h43a: dout <=  'sd2282; // 1082
        'h43b: dout <=  'sd189; // 1083
        'h43c: dout <=  'sd328; // 1084
        'h43d: dout <=  'sd330; // 1085
        'h43e: dout <= -'sd107; // 1086
        'h43f: dout <=  'sd634; // 1087
        'h440: dout <= -'sd1321; // 1088
        'h441: dout <= -'sd1049; // 1089
        'h442: dout <=  'sd1662; // 1090
        'h443: dout <= -'sd366; // 1091
        'h444: dout <= -'sd2046; // 1092
        'h445: dout <= -'sd772; // 1093
        'h446: dout <= -'sd1628; // 1094
        'h447: dout <= -'sd1301; // 1095
        'h448: dout <= -'sd116; // 1096
        'h449: dout <=  'sd139; // 1097
        'h44a: dout <=  'sd1003; // 1098
        'h44b: dout <=  'sd425; // 1099
        'h44c: dout <= -'sd901; // 1100
        'h44d: dout <=  'sd2248; // 1101
        'h44e: dout <= -'sd86; // 1102
        'h44f: dout <=  'sd62; // 1103
        'h450: dout <= -'sd1863; // 1104
        'h451: dout <= -'sd1533; // 1105
        'h452: dout <= -'sd245; // 1106
        'h453: dout <= -'sd321; // 1107
        'h454: dout <=  'sd1541; // 1108
        'h455: dout <= -'sd1040; // 1109
        'h456: dout <=  'sd2148; // 1110
        'h457: dout <= -'sd2021; // 1111
        'h458: dout <=  'sd104; // 1112
        'h459: dout <= -'sd2112; // 1113
        'h45a: dout <=  'sd1548; // 1114
        'h45b: dout <= -'sd796; // 1115
        'h45c: dout <= -'sd1468; // 1116
        'h45d: dout <= -'sd1621; // 1117
        'h45e: dout <= -'sd593; // 1118
        'h45f: dout <=  'sd343; // 1119
        'h460: dout <=  'sd263; // 1120
        'h461: dout <=  'sd1645; // 1121
        'h462: dout <= -'sd1289; // 1122
        'h463: dout <=  'sd2211; // 1123
        'h464: dout <=  'sd2281; // 1124
        'h465: dout <=  'sd684; // 1125
        'h466: dout <=  'sd1439; // 1126
        'h467: dout <=  'sd1106; // 1127
        'h468: dout <=  'sd1584; // 1128
        'h469: dout <=  'sd2094; // 1129
        'h46a: dout <=  'sd976; // 1130
        'h46b: dout <=  'sd1607; // 1131
        'h46c: dout <=  'sd2085; // 1132
        'h46d: dout <= -'sd1577; // 1133
        'h46e: dout <= -'sd2238; // 1134
        'h46f: dout <=  'sd1215; // 1135
        'h470: dout <=  'sd2292; // 1136
        'h471: dout <= -'sd14; // 1137
        'h472: dout <= -'sd1945; // 1138
        'h473: dout <=  'sd2072; // 1139
        'h474: dout <= -'sd840; // 1140
        'h475: dout <= -'sd349; // 1141
        'h476: dout <= -'sd646; // 1142
        'h477: dout <= -'sd1516; // 1143
        'h478: dout <= -'sd1634; // 1144
        'h479: dout <= -'sd575; // 1145
        'h47a: dout <=  'sd405; // 1146
        'h47b: dout <= -'sd1688; // 1147
        'h47c: dout <= -'sd1777; // 1148
        'h47d: dout <=  'sd433; // 1149
        'h47e: dout <=  'sd2237; // 1150
        'h47f: dout <= -'sd910; // 1151
        'h480: dout <=  'sd1007; // 1152
        'h481: dout <=  'sd852; // 1153
        'h482: dout <= -'sd2132; // 1154
        'h483: dout <=  'sd1338; // 1155
        'h484: dout <=  'sd1643; // 1156
        'h485: dout <=  'sd152; // 1157
        'h486: dout <=  'sd2183; // 1158
        'h487: dout <= -'sd1222; // 1159
        'h488: dout <= -'sd249; // 1160
        'h489: dout <= -'sd1438; // 1161
        'h48a: dout <=  'sd560; // 1162
        'h48b: dout <= -'sd908; // 1163
        'h48c: dout <= -'sd2178; // 1164
        'h48d: dout <=  'sd1838; // 1165
        'h48e: dout <= -'sd1755; // 1166
        'h48f: dout <= -'sd1682; // 1167
        'h490: dout <= -'sd1422; // 1168
        'h491: dout <=  'sd292; // 1169
        'h492: dout <= -'sd1250; // 1170
        'h493: dout <= -'sd1492; // 1171
        'h494: dout <= -'sd567; // 1172
        'h495: dout <= -'sd2049; // 1173
        'h496: dout <= -'sd1225; // 1174
        'h497: dout <=  'sd1175; // 1175
        'h498: dout <= -'sd1669; // 1176
        'h499: dout <= -'sd1610; // 1177
        'h49a: dout <=  'sd825; // 1178
        'h49b: dout <= -'sd2263; // 1179
        'h49c: dout <=  'sd359; // 1180
        'h49d: dout <=  'sd1569; // 1181
        'h49e: dout <=  'sd2079; // 1182
        'h49f: dout <=  'sd2059; // 1183
        'h4a0: dout <= -'sd1868; // 1184
        'h4a1: dout <=  'sd2002; // 1185
        'h4a2: dout <=  'sd1153; // 1186
        'h4a3: dout <=  'sd286; // 1187
        'h4a4: dout <= -'sd87; // 1188
        'h4a5: dout <= -'sd2163; // 1189
        'h4a6: dout <=  'sd2018; // 1190
        'h4a7: dout <=  'sd661; // 1191
        'h4a8: dout <=  'sd656; // 1192
        'h4a9: dout <=  'sd1525; // 1193
        'h4aa: dout <= -'sd1607; // 1194
        'h4ab: dout <=  'sd706; // 1195
        'h4ac: dout <= -'sd2243; // 1196
        'h4ad: dout <=  'sd899; // 1197
        'h4ae: dout <= -'sd1630; // 1198
        'h4af: dout <=  'sd1336; // 1199
        'h4b0: dout <= -'sd655; // 1200
        'h4b1: dout <=  'sd979; // 1201
        'h4b2: dout <=  'sd1976; // 1202
        'h4b3: dout <= -'sd644; // 1203
        'h4b4: dout <= -'sd787; // 1204
        'h4b5: dout <= -'sd2061; // 1205
        'h4b6: dout <= -'sd1214; // 1206
        'h4b7: dout <=  'sd471; // 1207
        'h4b8: dout <= -'sd1270; // 1208
        'h4b9: dout <=  'sd1533; // 1209
        'h4ba: dout <= -'sd53; // 1210
        'h4bb: dout <=  'sd267; // 1211
        'h4bc: dout <= -'sd284; // 1212
        'h4bd: dout <=  'sd243; // 1213
        'h4be: dout <= -'sd2023; // 1214
        'h4bf: dout <= -'sd928; // 1215
        'h4c0: dout <= -'sd1249; // 1216
        'h4c1: dout <=  'sd2197; // 1217
        'h4c2: dout <= -'sd360; // 1218
        'h4c3: dout <= -'sd1738; // 1219
        'h4c4: dout <=  'sd1914; // 1220
        'h4c5: dout <=  'sd1591; // 1221
        'h4c6: dout <= -'sd654; // 1222
        'h4c7: dout <=  'sd2185; // 1223
        'h4c8: dout <= -'sd78; // 1224
        'h4c9: dout <= -'sd804; // 1225
        'h4ca: dout <=  'sd1215; // 1226
        'h4cb: dout <= -'sd2127; // 1227
        'h4cc: dout <= -'sd399; // 1228
        'h4cd: dout <= -'sd1704; // 1229
        'h4ce: dout <=  'sd209; // 1230
        'h4cf: dout <=  'sd1155; // 1231
        'h4d0: dout <=  'sd1570; // 1232
        'h4d1: dout <= -'sd98; // 1233
        'h4d2: dout <=  'sd694; // 1234
        'h4d3: dout <=  'sd2283; // 1235
        'h4d4: dout <= -'sd218; // 1236
        'h4d5: dout <=  'sd1635; // 1237
        'h4d6: dout <= -'sd594; // 1238
        'h4d7: dout <=  'sd382; // 1239
        'h4d8: dout <= -'sd2050; // 1240
        'h4d9: dout <= -'sd2221; // 1241
        'h4da: dout <= -'sd1236; // 1242
        'h4db: dout <=  'sd160; // 1243
        'h4dc: dout <=  'sd1216; // 1244
        'h4dd: dout <=  'sd1577; // 1245
        'h4de: dout <=  'sd1792; // 1246
        'h4df: dout <= -'sd752; // 1247
        'h4e0: dout <= -'sd292; // 1248
        'h4e1: dout <= -'sd1708; // 1249
        'h4e2: dout <= -'sd1051; // 1250
        'h4e3: dout <=  'sd526; // 1251
        'h4e4: dout <=  'sd489; // 1252
        'h4e5: dout <= -'sd1552; // 1253
        'h4e6: dout <=  'sd355; // 1254
        'h4e7: dout <=  'sd1121; // 1255
        'h4e8: dout <= -'sd475; // 1256
        'h4e9: dout <= -'sd2217; // 1257
        'h4ea: dout <=  'sd1275; // 1258
        'h4eb: dout <=  'sd45; // 1259
        'h4ec: dout <= -'sd1977; // 1260
        'h4ed: dout <=  'sd419; // 1261
        'h4ee: dout <= -'sd63; // 1262
        'h4ef: dout <=  'sd1323; // 1263
        'h4f0: dout <=  'sd867; // 1264
        'h4f1: dout <= -'sd1527; // 1265
        'h4f2: dout <=  'sd1430; // 1266
        'h4f3: dout <= -'sd1790; // 1267
        'h4f4: dout <=  'sd18; // 1268
        'h4f5: dout <=  'sd1502; // 1269
        'h4f6: dout <= -'sd2038; // 1270
        'h4f7: dout <= -'sd1933; // 1271
        'h4f8: dout <= -'sd1423; // 1272
        'h4f9: dout <= -'sd927; // 1273
        'h4fa: dout <= -'sd22; // 1274
        'h4fb: dout <= -'sd1244; // 1275
        'h4fc: dout <=  'sd1771; // 1276
        'h4fd: dout <=  'sd1722; // 1277
        'h4fe: dout <= -'sd1321; // 1278
        'h4ff: dout <=  'sd1750; // 1279
        'h500: dout <=  'sd1917; // 1280
        'h501: dout <= -'sd1610; // 1281
        'h502: dout <= -'sd748; // 1282
        'h503: dout <=  'sd1600; // 1283
        'h504: dout <=  'sd1532; // 1284
        'h505: dout <= -'sd1269; // 1285
        'h506: dout <=  'sd1485; // 1286
        'h507: dout <= -'sd731; // 1287
        'h508: dout <= -'sd2014; // 1288
        'h509: dout <=  'sd454; // 1289
        'h50a: dout <=  'sd1054; // 1290
        'h50b: dout <=  'sd1492; // 1291
        'h50c: dout <= -'sd615; // 1292
        'h50d: dout <= -'sd1102; // 1293
        'h50e: dout <=  'sd2180; // 1294
        'h50f: dout <= -'sd1727; // 1295
        'h510: dout <=  'sd1192; // 1296
        'h511: dout <=  'sd797; // 1297
        'h512: dout <= -'sd513; // 1298
        'h513: dout <=  'sd675; // 1299
        'h514: dout <=  'sd1429; // 1300
        'h515: dout <=  'sd1624; // 1301
        'h516: dout <=  'sd745; // 1302
        'h517: dout <=  'sd1725; // 1303
        'h518: dout <= -'sd1010; // 1304
        'h519: dout <=  'sd302; // 1305
        'h51a: dout <=  'sd1733; // 1306
        'h51b: dout <=  'sd879; // 1307
        'h51c: dout <= -'sd925; // 1308
        'h51d: dout <= -'sd352; // 1309
        'h51e: dout <=  'sd916; // 1310
        'h51f: dout <= -'sd1260; // 1311
        'h520: dout <=  'sd1305; // 1312
        'h521: dout <=  'sd1384; // 1313
        'h522: dout <=  'sd2040; // 1314
        'h523: dout <= -'sd2271; // 1315
        'h524: dout <=  'sd944; // 1316
        'h525: dout <=  'sd652; // 1317
        'h526: dout <= -'sd1962; // 1318
        'h527: dout <=  'sd293; // 1319
        'h528: dout <=  'sd1637; // 1320
        'h529: dout <=  'sd1074; // 1321
        'h52a: dout <=  'sd1950; // 1322
        'h52b: dout <=  'sd1414; // 1323
        'h52c: dout <=  'sd205; // 1324
        'h52d: dout <= -'sd2012; // 1325
        'h52e: dout <=  'sd1811; // 1326
        'h52f: dout <= -'sd1270; // 1327
        'h530: dout <= -'sd947; // 1328
        'h531: dout <=  'sd1323; // 1329
        'h532: dout <= -'sd1962; // 1330
        'h533: dout <=  'sd171; // 1331
        'h534: dout <=  'sd984; // 1332
        'h535: dout <= -'sd1738; // 1333
        'h536: dout <= -'sd1009; // 1334
        'h537: dout <=  'sd1445; // 1335
        'h538: dout <=  'sd1657; // 1336
        'h539: dout <=  'sd1983; // 1337
        'h53a: dout <=  'sd1309; // 1338
        'h53b: dout <=  'sd1791; // 1339
        'h53c: dout <= -'sd2224; // 1340
        'h53d: dout <= -'sd2103; // 1341
        'h53e: dout <=  'sd1736; // 1342
        'h53f: dout <=  'sd1572; // 1343
        'h540: dout <= -'sd2071; // 1344
        'h541: dout <=  'sd1898; // 1345
        'h542: dout <=  'sd73; // 1346
        'h543: dout <=  'sd84; // 1347
        'h544: dout <=  'sd515; // 1348
        'h545: dout <=  'sd571; // 1349
        'h546: dout <= -'sd922; // 1350
        'h547: dout <=  'sd679; // 1351
        'h548: dout <= -'sd819; // 1352
        'h549: dout <= -'sd339; // 1353
        'h54a: dout <=  'sd2269; // 1354
        'h54b: dout <=  'sd598; // 1355
        'h54c: dout <=  'sd1983; // 1356
        'h54d: dout <= -'sd301; // 1357
        'h54e: dout <= -'sd1113; // 1358
        'h54f: dout <=  'sd329; // 1359
        'h550: dout <= -'sd1790; // 1360
        'h551: dout <= -'sd2246; // 1361
        'h552: dout <=  'sd1019; // 1362
        'h553: dout <= -'sd1043; // 1363
        'h554: dout <=  'sd1859; // 1364
        'h555: dout <=  'sd1139; // 1365
        'h556: dout <= -'sd1353; // 1366
        'h557: dout <=  'sd1062; // 1367
        'h558: dout <=  'sd1847; // 1368
        'h559: dout <= -'sd2224; // 1369
        'h55a: dout <= -'sd1882; // 1370
        'h55b: dout <= -'sd796; // 1371
        'h55c: dout <= -'sd1516; // 1372
        'h55d: dout <= -'sd2169; // 1373
        'h55e: dout <=  'sd2215; // 1374
        'h55f: dout <=  'sd341; // 1375
        'h560: dout <=  'sd952; // 1376
        'h561: dout <= -'sd1057; // 1377
        'h562: dout <= -'sd163; // 1378
        'h563: dout <= -'sd1067; // 1379
        'h564: dout <= -'sd2028; // 1380
        'h565: dout <=  'sd608; // 1381
        'h566: dout <=  'sd1440; // 1382
        'h567: dout <=  'sd1288; // 1383
        'h568: dout <= -'sd2050; // 1384
        'h569: dout <=  'sd2126; // 1385
        'h56a: dout <=  'sd80; // 1386
        'h56b: dout <=  'sd1055; // 1387
        'h56c: dout <=  'sd632; // 1388
        'h56d: dout <=  'sd1932; // 1389
        'h56e: dout <= -'sd505; // 1390
        'h56f: dout <= -'sd1622; // 1391
        'h570: dout <=  'sd1566; // 1392
        'h571: dout <= -'sd639; // 1393
        'h572: dout <=  'sd1219; // 1394
        'h573: dout <= -'sd188; // 1395
        'h574: dout <=  'sd647; // 1396
        'h575: dout <=  'sd601; // 1397
        'h576: dout <= -'sd966; // 1398
        'h577: dout <= -'sd670; // 1399
        'h578: dout <= -'sd1303; // 1400
        'h579: dout <= -'sd848; // 1401
        'h57a: dout <= -'sd1632; // 1402
        'h57b: dout <=  'sd2101; // 1403
        'h57c: dout <= -'sd1609; // 1404
        'h57d: dout <= -'sd414; // 1405
        'h57e: dout <= -'sd1278; // 1406
        'h57f: dout <= -'sd1102; // 1407
        'h580: dout <=  'sd1325; // 1408
        'h581: dout <=  'sd12; // 1409
        'h582: dout <= -'sd1393; // 1410
        'h583: dout <= -'sd1615; // 1411
        'h584: dout <=  'sd1077; // 1412
        'h585: dout <= -'sd376; // 1413
        'h586: dout <=  'sd1478; // 1414
        'h587: dout <=  'sd106; // 1415
        'h588: dout <= -'sd2063; // 1416
        'h589: dout <= -'sd1415; // 1417
        'h58a: dout <=  'sd1518; // 1418
        'h58b: dout <= -'sd1444; // 1419
        'h58c: dout <= -'sd1511; // 1420
        'h58d: dout <=  'sd1806; // 1421
        'h58e: dout <=  'sd1865; // 1422
        'h58f: dout <=  'sd1422; // 1423
        'h590: dout <=  'sd44; // 1424
        'h591: dout <= -'sd850; // 1425
        'h592: dout <=  'sd2159; // 1426
        'h593: dout <= -'sd920; // 1427
        'h594: dout <= -'sd257; // 1428
        'h595: dout <= -'sd1940; // 1429
        'h596: dout <= -'sd1254; // 1430
        'h597: dout <=  'sd823; // 1431
        'h598: dout <= -'sd152; // 1432
        'h599: dout <= -'sd720; // 1433
        'h59a: dout <=  'sd1429; // 1434
        'h59b: dout <=  'sd2023; // 1435
        'h59c: dout <=  'sd1483; // 1436
        'h59d: dout <=  'sd1885; // 1437
        'h59e: dout <=  'sd488; // 1438
        'h59f: dout <= -'sd305; // 1439
        'h5a0: dout <=  'sd684; // 1440
        'h5a1: dout <=  'sd370; // 1441
        'h5a2: dout <= -'sd894; // 1442
        'h5a3: dout <=  'sd1373; // 1443
        'h5a4: dout <= -'sd319; // 1444
        'h5a5: dout <= -'sd1866; // 1445
        'h5a6: dout <=  'sd897; // 1446
        'h5a7: dout <=  'sd1134; // 1447
        'h5a8: dout <= -'sd119; // 1448
        'h5a9: dout <=  'sd83; // 1449
        'h5aa: dout <=  'sd887; // 1450
        'h5ab: dout <=  'sd1696; // 1451
        'h5ac: dout <= -'sd851; // 1452
        'h5ad: dout <=  'sd1563; // 1453
        'h5ae: dout <=  'sd831; // 1454
        'h5af: dout <= -'sd518; // 1455
        'h5b0: dout <= -'sd474; // 1456
        'h5b1: dout <=  'sd210; // 1457
        'h5b2: dout <=  'sd582; // 1458
        'h5b3: dout <=  'sd4; // 1459
        'h5b4: dout <= -'sd1812; // 1460
        'h5b5: dout <= -'sd610; // 1461
        'h5b6: dout <= -'sd2258; // 1462
        'h5b7: dout <=  'sd137; // 1463
        'h5b8: dout <= -'sd1900; // 1464
        'h5b9: dout <=  'sd358; // 1465
        'h5ba: dout <=  'sd2136; // 1466
        'h5bb: dout <= -'sd345; // 1467
        'h5bc: dout <= -'sd135; // 1468
        'h5bd: dout <= -'sd297; // 1469
        'h5be: dout <=  'sd1242; // 1470
        'h5bf: dout <= -'sd179; // 1471
        'h5c0: dout <=  'sd812; // 1472
        'h5c1: dout <= -'sd1565; // 1473
        'h5c2: dout <=  'sd1983; // 1474
        'h5c3: dout <= -'sd881; // 1475
        'h5c4: dout <= -'sd2205; // 1476
        'h5c5: dout <= -'sd1107; // 1477
        'h5c6: dout <=  'sd460; // 1478
        'h5c7: dout <= -'sd2115; // 1479
        'h5c8: dout <= -'sd117; // 1480
        'h5c9: dout <= -'sd1128; // 1481
        'h5ca: dout <= -'sd1752; // 1482
        'h5cb: dout <=  'sd2205; // 1483
        'h5cc: dout <= -'sd2029; // 1484
        'h5cd: dout <= -'sd1112; // 1485
        'h5ce: dout <=  'sd1526; // 1486
        'h5cf: dout <=  'sd2178; // 1487
        'h5d0: dout <=  'sd7; // 1488
        'h5d1: dout <=  'sd1965; // 1489
        'h5d2: dout <= -'sd1513; // 1490
        'h5d3: dout <= -'sd725; // 1491
        'h5d4: dout <=  'sd1480; // 1492
        'h5d5: dout <= -'sd982; // 1493
        'h5d6: dout <=  'sd1661; // 1494
        'h5d7: dout <= -'sd2216; // 1495
        'h5d8: dout <= -'sd1819; // 1496
        'h5d9: dout <=  'sd165; // 1497
        'h5da: dout <=  'sd1427; // 1498
        'h5db: dout <= -'sd754; // 1499
        'h5dc: dout <= -'sd2227; // 1500
        'h5dd: dout <=  'sd901; // 1501
        'h5de: dout <=  'sd644; // 1502
        'h5df: dout <= -'sd277; // 1503
        'h5e0: dout <= -'sd1130; // 1504
        'h5e1: dout <= -'sd266; // 1505
        'h5e2: dout <= -'sd796; // 1506
        'h5e3: dout <=  'sd664; // 1507
        'h5e4: dout <= -'sd471; // 1508
        'h5e5: dout <= -'sd1280; // 1509
        'h5e6: dout <= -'sd2246; // 1510
        'h5e7: dout <= -'sd2033; // 1511
        'h5e8: dout <= -'sd1614; // 1512
        'h5e9: dout <= -'sd268; // 1513
        'h5ea: dout <=  'sd593; // 1514
        'h5eb: dout <=  'sd315; // 1515
        'h5ec: dout <=  'sd1994; // 1516
        'h5ed: dout <=  'sd1152; // 1517
        'h5ee: dout <=  'sd1485; // 1518
        'h5ef: dout <= -'sd2210; // 1519
        'h5f0: dout <=  'sd1335; // 1520
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hp_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [12:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <=  'sd727; // 0
        'h001: dout <=  'sd936; // 1
        'h002: dout <=  'sd1795; // 2
        'h003: dout <=  'sd48; // 3
        'h004: dout <= -'sd1549; // 4
        'h005: dout <= -'sd814; // 5
        'h006: dout <= -'sd1230; // 6
        'h007: dout <= -'sd1301; // 7
        'h008: dout <=  'sd1068; // 8
        'h009: dout <=  'sd471; // 9
        'h00a: dout <=  'sd314; // 10
        'h00b: dout <= -'sd383; // 11
        'h00c: dout <=  'sd1260; // 12
        'h00d: dout <= -'sd1382; // 13
        'h00e: dout <= -'sd1737; // 14
        'h00f: dout <= -'sd2049; // 15
        'h010: dout <= -'sd2192; // 16
        'h011: dout <= -'sd721; // 17
        'h012: dout <= -'sd1742; // 18
        'h013: dout <= -'sd1102; // 19
        'h014: dout <= -'sd508; // 20
        'h015: dout <= -'sd982; // 21
        'h016: dout <= -'sd733; // 22
        'h017: dout <= -'sd1626; // 23
        'h018: dout <= -'sd2236; // 24
        'h019: dout <= -'sd1070; // 25
        'h01a: dout <=  'sd1752; // 26
        'h01b: dout <=  'sd2280; // 27
        'h01c: dout <= -'sd1562; // 28
        'h01d: dout <=  'sd1866; // 29
        'h01e: dout <= -'sd1334; // 30
        'h01f: dout <= -'sd2199; // 31
        'h020: dout <=  'sd127; // 32
        'h021: dout <= -'sd89; // 33
        'h022: dout <= -'sd213; // 34
        'h023: dout <= -'sd432; // 35
        'h024: dout <=  'sd1921; // 36
        'h025: dout <= -'sd1002; // 37
        'h026: dout <=  'sd1726; // 38
        'h027: dout <= -'sd1803; // 39
        'h028: dout <=  'sd1049; // 40
        'h029: dout <=  'sd1464; // 41
        'h02a: dout <=  'sd1992; // 42
        'h02b: dout <= -'sd1499; // 43
        'h02c: dout <=  'sd1255; // 44
        'h02d: dout <=  'sd904; // 45
        'h02e: dout <= -'sd2069; // 46
        'h02f: dout <= -'sd842; // 47
        'h030: dout <= -'sd78; // 48
        'h031: dout <=  'sd931; // 49
        'h032: dout <= -'sd293; // 50
        'h033: dout <=  'sd1875; // 51
        'h034: dout <=  'sd1882; // 52
        'h035: dout <=  'sd1176; // 53
        'h036: dout <=  'sd1182; // 54
        'h037: dout <= -'sd389; // 55
        'h038: dout <= -'sd1232; // 56
        'h039: dout <= -'sd1605; // 57
        'h03a: dout <=  'sd1657; // 58
        'h03b: dout <=  'sd1421; // 59
        'h03c: dout <=  'sd139; // 60
        'h03d: dout <= -'sd247; // 61
        'h03e: dout <=  'sd828; // 62
        'h03f: dout <= -'sd850; // 63
        'h040: dout <=  'sd438; // 64
        'h041: dout <= -'sd456; // 65
        'h042: dout <=  'sd1197; // 66
        'h043: dout <=  'sd1082; // 67
        'h044: dout <=  'sd182; // 68
        'h045: dout <= -'sd2259; // 69
        'h046: dout <=  'sd851; // 70
        'h047: dout <=  'sd2245; // 71
        'h048: dout <= -'sd982; // 72
        'h049: dout <=  'sd139; // 73
        'h04a: dout <=  'sd827; // 74
        'h04b: dout <= -'sd1938; // 75
        'h04c: dout <= -'sd1297; // 76
        'h04d: dout <= -'sd1567; // 77
        'h04e: dout <= -'sd1708; // 78
        'h04f: dout <= -'sd534; // 79
        'h050: dout <=  'sd927; // 80
        'h051: dout <=  'sd845; // 81
        'h052: dout <= -'sd196; // 82
        'h053: dout <= -'sd1124; // 83
        'h054: dout <=  'sd1764; // 84
        'h055: dout <=  'sd1745; // 85
        'h056: dout <=  'sd324; // 86
        'h057: dout <= -'sd2120; // 87
        'h058: dout <= -'sd1069; // 88
        'h059: dout <= -'sd799; // 89
        'h05a: dout <=  'sd62; // 90
        'h05b: dout <= -'sd58; // 91
        'h05c: dout <=  'sd352; // 92
        'h05d: dout <= -'sd279; // 93
        'h05e: dout <=  'sd470; // 94
        'h05f: dout <=  'sd373; // 95
        'h060: dout <= -'sd317; // 96
        'h061: dout <= -'sd1328; // 97
        'h062: dout <=  'sd276; // 98
        'h063: dout <= -'sd648; // 99
        'h064: dout <=  'sd1313; // 100
        'h065: dout <=  'sd1216; // 101
        'h066: dout <= -'sd1247; // 102
        'h067: dout <= -'sd1629; // 103
        'h068: dout <= -'sd1055; // 104
        'h069: dout <=  'sd2145; // 105
        'h06a: dout <=  'sd619; // 106
        'h06b: dout <= -'sd2213; // 107
        'h06c: dout <=  'sd1039; // 108
        'h06d: dout <=  'sd534; // 109
        'h06e: dout <=  'sd49; // 110
        'h06f: dout <= -'sd1533; // 111
        'h070: dout <= -'sd1916; // 112
        'h071: dout <=  'sd28; // 113
        'h072: dout <= -'sd1978; // 114
        'h073: dout <= -'sd1544; // 115
        'h074: dout <=  'sd1781; // 116
        'h075: dout <= -'sd1546; // 117
        'h076: dout <= -'sd155; // 118
        'h077: dout <= -'sd1274; // 119
        'h078: dout <= -'sd1511; // 120
        'h079: dout <=  'sd1693; // 121
        'h07a: dout <=  'sd67; // 122
        'h07b: dout <= -'sd950; // 123
        'h07c: dout <=  'sd315; // 124
        'h07d: dout <=  'sd522; // 125
        'h07e: dout <= -'sd134; // 126
        'h07f: dout <= -'sd276; // 127
        'h080: dout <=  'sd1279; // 128
        'h081: dout <= -'sd1733; // 129
        'h082: dout <=  'sd1970; // 130
        'h083: dout <= -'sd1676; // 131
        'h084: dout <= -'sd1201; // 132
        'h085: dout <=  'sd1244; // 133
        'h086: dout <=  'sd379; // 134
        'h087: dout <=  'sd1746; // 135
        'h088: dout <=  'sd1278; // 136
        'h089: dout <=  'sd993; // 137
        'h08a: dout <= -'sd1091; // 138
        'h08b: dout <= -'sd1629; // 139
        'h08c: dout <=  'sd1010; // 140
        'h08d: dout <= -'sd1541; // 141
        'h08e: dout <= -'sd471; // 142
        'h08f: dout <= -'sd1757; // 143
        'h090: dout <= -'sd163; // 144
        'h091: dout <=  'sd1892; // 145
        'h092: dout <= -'sd938; // 146
        'h093: dout <= -'sd1447; // 147
        'h094: dout <= -'sd1710; // 148
        'h095: dout <= -'sd1730; // 149
        'h096: dout <=  'sd1732; // 150
        'h097: dout <= -'sd1352; // 151
        'h098: dout <=  'sd1227; // 152
        'h099: dout <= -'sd1022; // 153
        'h09a: dout <= -'sd667; // 154
        'h09b: dout <= -'sd467; // 155
        'h09c: dout <= -'sd282; // 156
        'h09d: dout <= -'sd2164; // 157
        'h09e: dout <= -'sd1994; // 158
        'h09f: dout <= -'sd1691; // 159
        'h0a0: dout <=  'sd997; // 160
        'h0a1: dout <= -'sd498; // 161
        'h0a2: dout <= -'sd366; // 162
        'h0a3: dout <= -'sd1607; // 163
        'h0a4: dout <= -'sd1719; // 164
        'h0a5: dout <=  'sd1486; // 165
        'h0a6: dout <=  'sd1328; // 166
        'h0a7: dout <= -'sd1841; // 167
        'h0a8: dout <=  'sd1004; // 168
        'h0a9: dout <=  'sd162; // 169
        'h0aa: dout <= -'sd1302; // 170
        'h0ab: dout <=  'sd762; // 171
        'h0ac: dout <= -'sd1038; // 172
        'h0ad: dout <= -'sd636; // 173
        'h0ae: dout <=  'sd2150; // 174
        'h0af: dout <= -'sd1612; // 175
        'h0b0: dout <=  'sd1191; // 176
        'h0b1: dout <=  'sd305; // 177
        'h0b2: dout <=  'sd1349; // 178
        'h0b3: dout <= -'sd330; // 179
        'h0b4: dout <=  'sd1057; // 180
        'h0b5: dout <=  'sd1207; // 181
        'h0b6: dout <= -'sd350; // 182
        'h0b7: dout <= -'sd676; // 183
        'h0b8: dout <=  'sd1217; // 184
        'h0b9: dout <=  'sd21; // 185
        'h0ba: dout <=  'sd199; // 186
        'h0bb: dout <= -'sd817; // 187
        'h0bc: dout <= -'sd966; // 188
        'h0bd: dout <=  'sd960; // 189
        'h0be: dout <= -'sd1186; // 190
        'h0bf: dout <=  'sd596; // 191
        'h0c0: dout <= -'sd918; // 192
        'h0c1: dout <=  'sd1229; // 193
        'h0c2: dout <=  'sd402; // 194
        'h0c3: dout <=  'sd165; // 195
        'h0c4: dout <= -'sd1446; // 196
        'h0c5: dout <=  'sd1450; // 197
        'h0c6: dout <= -'sd1572; // 198
        'h0c7: dout <=  'sd588; // 199
        'h0c8: dout <= -'sd2175; // 200
        'h0c9: dout <=  'sd54; // 201
        'h0ca: dout <=  'sd1827; // 202
        'h0cb: dout <= -'sd1884; // 203
        'h0cc: dout <= -'sd2146; // 204
        'h0cd: dout <=  'sd79; // 205
        'h0ce: dout <= -'sd1861; // 206
        'h0cf: dout <= -'sd515; // 207
        'h0d0: dout <= -'sd1665; // 208
        'h0d1: dout <= -'sd1857; // 209
        'h0d2: dout <= -'sd1391; // 210
        'h0d3: dout <= -'sd1631; // 211
        'h0d4: dout <=  'sd1020; // 212
        'h0d5: dout <= -'sd1387; // 213
        'h0d6: dout <= -'sd808; // 214
        'h0d7: dout <=  'sd560; // 215
        'h0d8: dout <= -'sd1448; // 216
        'h0d9: dout <=  'sd559; // 217
        'h0da: dout <= -'sd2178; // 218
        'h0db: dout <=  'sd673; // 219
        'h0dc: dout <= -'sd2063; // 220
        'h0dd: dout <= -'sd147; // 221
        'h0de: dout <= -'sd535; // 222
        'h0df: dout <= -'sd427; // 223
        'h0e0: dout <= -'sd633; // 224
        'h0e1: dout <= -'sd705; // 225
        'h0e2: dout <= -'sd1882; // 226
        'h0e3: dout <=  'sd662; // 227
        'h0e4: dout <=  'sd531; // 228
        'h0e5: dout <=  'sd1280; // 229
        'h0e6: dout <= -'sd409; // 230
        'h0e7: dout <=  'sd1009; // 231
        'h0e8: dout <=  'sd447; // 232
        'h0e9: dout <= -'sd2092; // 233
        'h0ea: dout <=  'sd2064; // 234
        'h0eb: dout <= -'sd13; // 235
        'h0ec: dout <= -'sd1457; // 236
        'h0ed: dout <=  'sd1575; // 237
        'h0ee: dout <=  'sd1525; // 238
        'h0ef: dout <= -'sd2243; // 239
        'h0f0: dout <= -'sd613; // 240
        'h0f1: dout <= -'sd117; // 241
        'h0f2: dout <=  'sd1258; // 242
        'h0f3: dout <= -'sd1868; // 243
        'h0f4: dout <=  'sd2198; // 244
        'h0f5: dout <= -'sd1977; // 245
        'h0f6: dout <= -'sd1308; // 246
        'h0f7: dout <=  'sd1762; // 247
        'h0f8: dout <=  'sd509; // 248
        'h0f9: dout <=  'sd1899; // 249
        'h0fa: dout <=  'sd1677; // 250
        'h0fb: dout <=  'sd357; // 251
        'h0fc: dout <= -'sd2221; // 252
        'h0fd: dout <= -'sd451; // 253
        'h0fe: dout <= -'sd339; // 254
        'h0ff: dout <= -'sd2171; // 255
        'h100: dout <=  'sd1895; // 256
        'h101: dout <= -'sd282; // 257
        'h102: dout <= -'sd630; // 258
        'h103: dout <=  'sd704; // 259
        'h104: dout <= -'sd1228; // 260
        'h105: dout <=  'sd1934; // 261
        'h106: dout <=  'sd807; // 262
        'h107: dout <=  'sd2158; // 263
        'h108: dout <= -'sd1991; // 264
        'h109: dout <=  'sd1814; // 265
        'h10a: dout <= -'sd2053; // 266
        'h10b: dout <=  'sd780; // 267
        'h10c: dout <=  'sd1315; // 268
        'h10d: dout <= -'sd964; // 269
        'h10e: dout <= -'sd1254; // 270
        'h10f: dout <= -'sd1049; // 271
        'h110: dout <= -'sd1006; // 272
        'h111: dout <= -'sd2246; // 273
        'h112: dout <= -'sd957; // 274
        'h113: dout <= -'sd1422; // 275
        'h114: dout <=  'sd1597; // 276
        'h115: dout <=  'sd674; // 277
        'h116: dout <= -'sd646; // 278
        'h117: dout <=  'sd137; // 279
        'h118: dout <= -'sd1542; // 280
        'h119: dout <= -'sd1048; // 281
        'h11a: dout <=  'sd220; // 282
        'h11b: dout <= -'sd564; // 283
        'h11c: dout <=  'sd709; // 284
        'h11d: dout <=  'sd1456; // 285
        'h11e: dout <=  'sd1480; // 286
        'h11f: dout <=  'sd7; // 287
        'h120: dout <=  'sd828; // 288
        'h121: dout <=  'sd1844; // 289
        'h122: dout <=  'sd1382; // 290
        'h123: dout <= -'sd351; // 291
        'h124: dout <=  'sd575; // 292
        'h125: dout <=  'sd429; // 293
        'h126: dout <= -'sd761; // 294
        'h127: dout <=  'sd239; // 295
        'h128: dout <= -'sd2069; // 296
        'h129: dout <= -'sd1729; // 297
        'h12a: dout <=  'sd1127; // 298
        'h12b: dout <= -'sd1889; // 299
        'h12c: dout <=  'sd854; // 300
        'h12d: dout <= -'sd743; // 301
        'h12e: dout <=  'sd1750; // 302
        'h12f: dout <= -'sd1899; // 303
        'h130: dout <=  'sd2284; // 304
        'h131: dout <=  'sd233; // 305
        'h132: dout <= -'sd398; // 306
        'h133: dout <= -'sd561; // 307
        'h134: dout <=  'sd215; // 308
        'h135: dout <= -'sd59; // 309
        'h136: dout <=  'sd1372; // 310
        'h137: dout <= -'sd552; // 311
        'h138: dout <=  'sd2128; // 312
        'h139: dout <=  'sd73; // 313
        'h13a: dout <= -'sd1825; // 314
        'h13b: dout <=  'sd616; // 315
        'h13c: dout <= -'sd1680; // 316
        'h13d: dout <=  'sd1338; // 317
        'h13e: dout <= -'sd389; // 318
        'h13f: dout <=  'sd402; // 319
        'h140: dout <=  'sd1222; // 320
        'h141: dout <= -'sd1977; // 321
        'h142: dout <=  'sd747; // 322
        'h143: dout <= -'sd1566; // 323
        'h144: dout <=  'sd1533; // 324
        'h145: dout <=  'sd2083; // 325
        'h146: dout <= -'sd1170; // 326
        'h147: dout <=  'sd786; // 327
        'h148: dout <= -'sd2263; // 328
        'h149: dout <= -'sd1535; // 329
        'h14a: dout <= -'sd977; // 330
        'h14b: dout <= -'sd208; // 331
        'h14c: dout <=  'sd2108; // 332
        'h14d: dout <= -'sd1693; // 333
        'h14e: dout <=  'sd1620; // 334
        'h14f: dout <= -'sd1978; // 335
        'h150: dout <=  'sd2267; // 336
        'h151: dout <= -'sd1983; // 337
        'h152: dout <= -'sd1590; // 338
        'h153: dout <= -'sd2243; // 339
        'h154: dout <= -'sd803; // 340
        'h155: dout <= -'sd1013; // 341
        'h156: dout <= -'sd2056; // 342
        'h157: dout <=  'sd1671; // 343
        'h158: dout <= -'sd1572; // 344
        'h159: dout <= -'sd2131; // 345
        'h15a: dout <=  'sd1424; // 346
        'h15b: dout <=  'sd1172; // 347
        'h15c: dout <=  'sd1244; // 348
        'h15d: dout <=  'sd2197; // 349
        'h15e: dout <=  'sd2109; // 350
        'h15f: dout <= -'sd87; // 351
        'h160: dout <=  'sd1050; // 352
        'h161: dout <=  'sd1493; // 353
        'h162: dout <=  'sd1791; // 354
        'h163: dout <= -'sd1897; // 355
        'h164: dout <= -'sd727; // 356
        'h165: dout <= -'sd1563; // 357
        'h166: dout <= -'sd1743; // 358
        'h167: dout <=  'sd2065; // 359
        'h168: dout <= -'sd1992; // 360
        'h169: dout <= -'sd505; // 361
        'h16a: dout <= -'sd1467; // 362
        'h16b: dout <= -'sd718; // 363
        'h16c: dout <= -'sd822; // 364
        'h16d: dout <= -'sd541; // 365
        'h16e: dout <=  'sd342; // 366
        'h16f: dout <=  'sd238; // 367
        'h170: dout <=  'sd2252; // 368
        'h171: dout <=  'sd1017; // 369
        'h172: dout <=  'sd367; // 370
        'h173: dout <=  'sd175; // 371
        'h174: dout <=  'sd1515; // 372
        'h175: dout <= -'sd2235; // 373
        'h176: dout <=  'sd1011; // 374
        'h177: dout <= -'sd1260; // 375
        'h178: dout <=  'sd466; // 376
        'h179: dout <=  'sd192; // 377
        'h17a: dout <=  'sd1901; // 378
        'h17b: dout <= -'sd840; // 379
        'h17c: dout <=  'sd343; // 380
        'h17d: dout <=  'sd1276; // 381
        'h17e: dout <=  'sd1434; // 382
        'h17f: dout <=  'sd1469; // 383
        'h180: dout <= -'sd326; // 384
        'h181: dout <=  'sd53; // 385
        'h182: dout <= -'sd1473; // 386
        'h183: dout <=  'sd1840; // 387
        'h184: dout <=  'sd708; // 388
        'h185: dout <=  'sd1839; // 389
        'h186: dout <=  'sd1943; // 390
        'h187: dout <=  'sd1886; // 391
        'h188: dout <= -'sd1516; // 392
        'h189: dout <=  'sd448; // 393
        'h18a: dout <=  'sd1129; // 394
        'h18b: dout <= -'sd1163; // 395
        'h18c: dout <=  'sd1349; // 396
        'h18d: dout <= -'sd15; // 397
        'h18e: dout <=  'sd396; // 398
        'h18f: dout <=  'sd1664; // 399
        'h190: dout <=  'sd1106; // 400
        'h191: dout <= -'sd1724; // 401
        'h192: dout <=  'sd751; // 402
        'h193: dout <=  'sd1552; // 403
        'h194: dout <=  'sd797; // 404
        'h195: dout <= -'sd399; // 405
        'h196: dout <=  'sd1191; // 406
        'h197: dout <= -'sd1852; // 407
        'h198: dout <=  'sd541; // 408
        'h199: dout <=  'sd359; // 409
        'h19a: dout <= -'sd2067; // 410
        'h19b: dout <= -'sd2059; // 411
        'h19c: dout <=  'sd1421; // 412
        'h19d: dout <=  'sd334; // 413
        'h19e: dout <= -'sd889; // 414
        'h19f: dout <=  'sd2038; // 415
        'h1a0: dout <=  'sd1113; // 416
        'h1a1: dout <=  'sd246; // 417
        'h1a2: dout <= -'sd412; // 418
        'h1a3: dout <= -'sd2212; // 419
        'h1a4: dout <=  'sd1742; // 420
        'h1a5: dout <= -'sd2214; // 421
        'h1a6: dout <= -'sd831; // 422
        'h1a7: dout <= -'sd2272; // 423
        'h1a8: dout <= -'sd465; // 424
        'h1a9: dout <= -'sd119; // 425
        'h1aa: dout <=  'sd2158; // 426
        'h1ab: dout <= -'sd25; // 427
        'h1ac: dout <=  'sd578; // 428
        'h1ad: dout <= -'sd1523; // 429
        'h1ae: dout <=  'sd1233; // 430
        'h1af: dout <= -'sd431; // 431
        'h1b0: dout <=  'sd882; // 432
        'h1b1: dout <= -'sd347; // 433
        'h1b2: dout <=  'sd1295; // 434
        'h1b3: dout <=  'sd1203; // 435
        'h1b4: dout <=  'sd989; // 436
        'h1b5: dout <=  'sd509; // 437
        'h1b6: dout <= -'sd515; // 438
        'h1b7: dout <= -'sd782; // 439
        'h1b8: dout <=  'sd808; // 440
        'h1b9: dout <= -'sd894; // 441
        'h1ba: dout <=  'sd815; // 442
        'h1bb: dout <=  'sd962; // 443
        'h1bc: dout <=  'sd1341; // 444
        'h1bd: dout <=  'sd80; // 445
        'h1be: dout <= -'sd2070; // 446
        'h1bf: dout <=  'sd1943; // 447
        'h1c0: dout <= -'sd1350; // 448
        'h1c1: dout <=  'sd112; // 449
        'h1c2: dout <= -'sd977; // 450
        'h1c3: dout <=  'sd385; // 451
        'h1c4: dout <=  'sd291; // 452
        'h1c5: dout <=  'sd1973; // 453
        'h1c6: dout <= -'sd308; // 454
        'h1c7: dout <=  'sd1590; // 455
        'h1c8: dout <= -'sd939; // 456
        'h1c9: dout <= -'sd1285; // 457
        'h1ca: dout <=  'sd543; // 458
        'h1cb: dout <=  'sd1329; // 459
        'h1cc: dout <=  'sd132; // 460
        'h1cd: dout <= -'sd425; // 461
        'h1ce: dout <=  'sd1554; // 462
        'h1cf: dout <=  'sd737; // 463
        'h1d0: dout <= -'sd740; // 464
        'h1d1: dout <=  'sd871; // 465
        'h1d2: dout <= -'sd2052; // 466
        'h1d3: dout <=  'sd574; // 467
        'h1d4: dout <=  'sd1998; // 468
        'h1d5: dout <=  'sd726; // 469
        'h1d6: dout <= -'sd74; // 470
        'h1d7: dout <= -'sd675; // 471
        'h1d8: dout <= -'sd820; // 472
        'h1d9: dout <=  'sd1744; // 473
        'h1da: dout <= -'sd1236; // 474
        'h1db: dout <=  'sd49; // 475
        'h1dc: dout <= -'sd1223; // 476
        'h1dd: dout <=  'sd1044; // 477
        'h1de: dout <=  'sd1066; // 478
        'h1df: dout <= -'sd1688; // 479
        'h1e0: dout <= -'sd1523; // 480
        'h1e1: dout <= -'sd1223; // 481
        'h1e2: dout <= -'sd800; // 482
        'h1e3: dout <= -'sd1476; // 483
        'h1e4: dout <=  'sd898; // 484
        'h1e5: dout <= -'sd1193; // 485
        'h1e6: dout <= -'sd1310; // 486
        'h1e7: dout <= -'sd578; // 487
        'h1e8: dout <= -'sd1692; // 488
        'h1e9: dout <= -'sd2188; // 489
        'h1ea: dout <=  'sd87; // 490
        'h1eb: dout <= -'sd2081; // 491
        'h1ec: dout <= -'sd1769; // 492
        'h1ed: dout <=  'sd1368; // 493
        'h1ee: dout <=  'sd263; // 494
        'h1ef: dout <=  'sd1250; // 495
        'h1f0: dout <=  'sd1808; // 496
        'h1f1: dout <=  'sd1356; // 497
        'h1f2: dout <=  'sd930; // 498
        'h1f3: dout <= -'sd1558; // 499
        'h1f4: dout <= -'sd2249; // 500
        'h1f5: dout <= -'sd2089; // 501
        'h1f6: dout <= -'sd82; // 502
        'h1f7: dout <=  'sd1320; // 503
        'h1f8: dout <= -'sd875; // 504
        'h1f9: dout <= -'sd2139; // 505
        'h1fa: dout <= -'sd810; // 506
        'h1fb: dout <=  'sd559; // 507
        'h1fc: dout <=  'sd2149; // 508
        'h1fd: dout <=  'sd2268; // 509
        'h1fe: dout <= -'sd1446; // 510
        'h1ff: dout <= -'sd1753; // 511
        'h200: dout <= -'sd1300; // 512
        'h201: dout <=  'sd2263; // 513
        'h202: dout <=  'sd127; // 514
        'h203: dout <=  'sd917; // 515
        'h204: dout <= -'sd16; // 516
        'h205: dout <=  'sd889; // 517
        'h206: dout <=  'sd1321; // 518
        'h207: dout <= -'sd1087; // 519
        'h208: dout <=  'sd617; // 520
        'h209: dout <= -'sd976; // 521
        'h20a: dout <=  'sd956; // 522
        'h20b: dout <= -'sd763; // 523
        'h20c: dout <= -'sd2287; // 524
        'h20d: dout <=  'sd59; // 525
        'h20e: dout <=  'sd1321; // 526
        'h20f: dout <=  'sd2035; // 527
        'h210: dout <= -'sd1292; // 528
        'h211: dout <=  'sd360; // 529
        'h212: dout <= -'sd1735; // 530
        'h213: dout <=  'sd117; // 531
        'h214: dout <=  'sd334; // 532
        'h215: dout <=  'sd1542; // 533
        'h216: dout <=  'sd1430; // 534
        'h217: dout <= -'sd1829; // 535
        'h218: dout <= -'sd1229; // 536
        'h219: dout <= -'sd853; // 537
        'h21a: dout <= -'sd1016; // 538
        'h21b: dout <= -'sd73; // 539
        'h21c: dout <=  'sd690; // 540
        'h21d: dout <= -'sd445; // 541
        'h21e: dout <=  'sd1002; // 542
        'h21f: dout <=  'sd1939; // 543
        'h220: dout <=  'sd453; // 544
        'h221: dout <=  'sd945; // 545
        'h222: dout <=  'sd1543; // 546
        'h223: dout <=  'sd192; // 547
        'h224: dout <= -'sd2253; // 548
        'h225: dout <=  'sd2219; // 549
        'h226: dout <= -'sd139; // 550
        'h227: dout <=  'sd2034; // 551
        'h228: dout <=  'sd839; // 552
        'h229: dout <= -'sd1984; // 553
        'h22a: dout <=  'sd244; // 554
        'h22b: dout <= -'sd5; // 555
        'h22c: dout <=  'sd2192; // 556
        'h22d: dout <=  'sd660; // 557
        'h22e: dout <= -'sd2093; // 558
        'h22f: dout <= -'sd2252; // 559
        'h230: dout <=  'sd2064; // 560
        'h231: dout <= -'sd626; // 561
        'h232: dout <=  'sd1175; // 562
        'h233: dout <= -'sd2289; // 563
        'h234: dout <=  'sd73; // 564
        'h235: dout <= -'sd291; // 565
        'h236: dout <=  'sd1748; // 566
        'h237: dout <=  'sd1356; // 567
        'h238: dout <= -'sd1848; // 568
        'h239: dout <= -'sd128; // 569
        'h23a: dout <= -'sd1849; // 570
        'h23b: dout <=  'sd278; // 571
        'h23c: dout <=  'sd1800; // 572
        'h23d: dout <=  'sd358; // 573
        'h23e: dout <=  'sd2175; // 574
        'h23f: dout <= -'sd1330; // 575
        'h240: dout <= -'sd1922; // 576
        'h241: dout <=  'sd549; // 577
        'h242: dout <= -'sd1412; // 578
        'h243: dout <= -'sd1574; // 579
        'h244: dout <= -'sd1032; // 580
        'h245: dout <= -'sd396; // 581
        'h246: dout <= -'sd1995; // 582
        'h247: dout <= -'sd644; // 583
        'h248: dout <= -'sd88; // 584
        'h249: dout <=  'sd1026; // 585
        'h24a: dout <=  'sd555; // 586
        'h24b: dout <=  'sd1261; // 587
        'h24c: dout <=  'sd343; // 588
        'h24d: dout <=  'sd309; // 589
        'h24e: dout <= -'sd462; // 590
        'h24f: dout <= -'sd1022; // 591
        'h250: dout <=  'sd1849; // 592
        'h251: dout <= -'sd1529; // 593
        'h252: dout <= -'sd2285; // 594
        'h253: dout <=  'sd2047; // 595
        'h254: dout <=  'sd935; // 596
        'h255: dout <=  'sd1914; // 597
        'h256: dout <= -'sd1151; // 598
        'h257: dout <=  'sd169; // 599
        'h258: dout <=  'sd945; // 600
        'h259: dout <=  'sd49; // 601
        'h25a: dout <=  'sd1691; // 602
        'h25b: dout <= -'sd1154; // 603
        'h25c: dout <= -'sd1513; // 604
        'h25d: dout <= -'sd2127; // 605
        'h25e: dout <= -'sd272; // 606
        'h25f: dout <=  'sd462; // 607
        'h260: dout <= -'sd2187; // 608
        'h261: dout <= -'sd756; // 609
        'h262: dout <= -'sd332; // 610
        'h263: dout <= -'sd1664; // 611
        'h264: dout <=  'sd1380; // 612
        'h265: dout <=  'sd1736; // 613
        'h266: dout <=  'sd1874; // 614
        'h267: dout <= -'sd764; // 615
        'h268: dout <= -'sd1316; // 616
        'h269: dout <= -'sd687; // 617
        'h26a: dout <=  'sd741; // 618
        'h26b: dout <= -'sd2200; // 619
        'h26c: dout <=  'sd1902; // 620
        'h26d: dout <=  'sd1434; // 621
        'h26e: dout <=  'sd175; // 622
        'h26f: dout <=  'sd2077; // 623
        'h270: dout <= -'sd206; // 624
        'h271: dout <=  'sd1322; // 625
        'h272: dout <= -'sd554; // 626
        'h273: dout <=  'sd395; // 627
        'h274: dout <=  'sd1763; // 628
        'h275: dout <= -'sd1635; // 629
        'h276: dout <=  'sd1978; // 630
        'h277: dout <= -'sd2046; // 631
        'h278: dout <=  'sd1968; // 632
        'h279: dout <=  'sd775; // 633
        'h27a: dout <=  'sd1916; // 634
        'h27b: dout <=  'sd564; // 635
        'h27c: dout <=  'sd112; // 636
        'h27d: dout <= -'sd178; // 637
        'h27e: dout <= -'sd1241; // 638
        'h27f: dout <= -'sd1975; // 639
        'h280: dout <=  'sd1572; // 640
        'h281: dout <=  'sd657; // 641
        'h282: dout <=  'sd519; // 642
        'h283: dout <= -'sd339; // 643
        'h284: dout <= -'sd295; // 644
        'h285: dout <=  'sd1483; // 645
        'h286: dout <=  'sd991; // 646
        'h287: dout <= -'sd2047; // 647
        'h288: dout <= -'sd1721; // 648
        'h289: dout <= -'sd125; // 649
        'h28a: dout <=  'sd1580; // 650
        'h28b: dout <= -'sd474; // 651
        'h28c: dout <=  'sd229; // 652
        'h28d: dout <=  'sd1724; // 653
        'h28e: dout <=  'sd1352; // 654
        'h28f: dout <= -'sd2021; // 655
        'h290: dout <= -'sd1061; // 656
        'h291: dout <= -'sd717; // 657
        'h292: dout <= -'sd110; // 658
        'h293: dout <= -'sd649; // 659
        'h294: dout <=  'sd1012; // 660
        'h295: dout <= -'sd567; // 661
        'h296: dout <=  'sd799; // 662
        'h297: dout <=  'sd1694; // 663
        'h298: dout <= -'sd334; // 664
        'h299: dout <=  'sd611; // 665
        'h29a: dout <=  'sd290; // 666
        'h29b: dout <= -'sd816; // 667
        'h29c: dout <= -'sd1101; // 668
        'h29d: dout <= -'sd2034; // 669
        'h29e: dout <=  'sd1680; // 670
        'h29f: dout <=  'sd673; // 671
        'h2a0: dout <=  'sd748; // 672
        'h2a1: dout <=  'sd1750; // 673
        'h2a2: dout <=  'sd174; // 674
        'h2a3: dout <= -'sd1291; // 675
        'h2a4: dout <= -'sd1880; // 676
        'h2a5: dout <=  'sd229; // 677
        'h2a6: dout <= -'sd1988; // 678
        'h2a7: dout <= -'sd917; // 679
        'h2a8: dout <= -'sd435; // 680
        'h2a9: dout <= -'sd1679; // 681
        'h2aa: dout <= -'sd170; // 682
        'h2ab: dout <= -'sd2229; // 683
        'h2ac: dout <=  'sd317; // 684
        'h2ad: dout <= -'sd494; // 685
        'h2ae: dout <=  'sd2268; // 686
        'h2af: dout <= -'sd109; // 687
        'h2b0: dout <= -'sd910; // 688
        'h2b1: dout <=  'sd1017; // 689
        'h2b2: dout <=  'sd2082; // 690
        'h2b3: dout <= -'sd1165; // 691
        'h2b4: dout <=  'sd650; // 692
        'h2b5: dout <=  'sd932; // 693
        'h2b6: dout <=  'sd518; // 694
        'h2b7: dout <= -'sd1097; // 695
        'h2b8: dout <= -'sd1095; // 696
        'h2b9: dout <= -'sd1647; // 697
        'h2ba: dout <= -'sd1241; // 698
        'h2bb: dout <=  'sd1713; // 699
        'h2bc: dout <= -'sd642; // 700
        'h2bd: dout <=  'sd2015; // 701
        'h2be: dout <= -'sd498; // 702
        'h2bf: dout <=  'sd768; // 703
        'h2c0: dout <= -'sd2258; // 704
        'h2c1: dout <= -'sd1893; // 705
        'h2c2: dout <= -'sd2082; // 706
        'h2c3: dout <=  'sd352; // 707
        'h2c4: dout <=  'sd1292; // 708
        'h2c5: dout <=  'sd1044; // 709
        'h2c6: dout <= -'sd1715; // 710
        'h2c7: dout <= -'sd291; // 711
        'h2c8: dout <= -'sd1968; // 712
        'h2c9: dout <= -'sd1895; // 713
        'h2ca: dout <=  'sd1017; // 714
        'h2cb: dout <=  'sd714; // 715
        'h2cc: dout <= -'sd1032; // 716
        'h2cd: dout <=  'sd385; // 717
        'h2ce: dout <=  'sd25; // 718
        'h2cf: dout <=  'sd2219; // 719
        'h2d0: dout <= -'sd695; // 720
        'h2d1: dout <=  'sd103; // 721
        'h2d2: dout <= -'sd1035; // 722
        'h2d3: dout <=  'sd1181; // 723
        'h2d4: dout <=  'sd1178; // 724
        'h2d5: dout <=  'sd1095; // 725
        'h2d6: dout <= -'sd1089; // 726
        'h2d7: dout <=  'sd518; // 727
        'h2d8: dout <= -'sd759; // 728
        'h2d9: dout <=  'sd1001; // 729
        'h2da: dout <= -'sd970; // 730
        'h2db: dout <=  'sd2113; // 731
        'h2dc: dout <= -'sd568; // 732
        'h2dd: dout <=  'sd811; // 733
        'h2de: dout <=  'sd1998; // 734
        'h2df: dout <= -'sd254; // 735
        'h2e0: dout <=  'sd575; // 736
        'h2e1: dout <=  'sd37; // 737
        'h2e2: dout <= -'sd233; // 738
        'h2e3: dout <=  'sd1669; // 739
        'h2e4: dout <=  'sd113; // 740
        'h2e5: dout <= -'sd128; // 741
        'h2e6: dout <=  'sd338; // 742
        'h2e7: dout <=  'sd2124; // 743
        'h2e8: dout <=  'sd572; // 744
        'h2e9: dout <=  'sd2013; // 745
        'h2ea: dout <=  'sd369; // 746
        'h2eb: dout <= -'sd703; // 747
        'h2ec: dout <=  'sd131; // 748
        'h2ed: dout <=  'sd773; // 749
        'h2ee: dout <=  'sd2110; // 750
        'h2ef: dout <= -'sd738; // 751
        'h2f0: dout <= -'sd1988; // 752
        'h2f1: dout <=  'sd1394; // 753
        'h2f2: dout <=  'sd2135; // 754
        'h2f3: dout <= -'sd2046; // 755
        'h2f4: dout <= -'sd98; // 756
        'h2f5: dout <=  'sd166; // 757
        'h2f6: dout <= -'sd876; // 758
        'h2f7: dout <= -'sd1869; // 759
        'h2f8: dout <= -'sd1044; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

