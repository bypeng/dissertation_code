module mod4591Svec33 (
    input       [32:0] z_in,
    output      [11:0] p0,
    output reg  [11:0] p1,
    output reg  [11:0] n0,
    output reg  [12:0] n1,
    output reg  [11:0] n2,
    output reg  [12:0] n3
) ;

    assign p0 = z_in[11:0];

    always @ (*) begin
        case({ z_in[32], z_in[23], z_in[18], z_in[15] })
            4'h0: p1 = 12'd0;
            4'h1: p1 = 12'd631;
            4'h2: p1 = 12'd457;
            4'h3: p1 = 12'd1088;
            4'h4: p1 = 12'd851;
            4'h5: p1 = 12'd1482;
            4'h6: p1 = 12'd1308;
            4'h7: p1 = 12'd1939;
            4'h8: p1 = 12'd433;
            4'h9: p1 = 12'd1064;
            4'ha: p1 = 12'd890;
            4'hb: p1 = 12'd1521;
            4'hc: p1 = 12'd1284;
            4'hd: p1 = 12'd1915;
            4'he: p1 = 12'd1741;
            4'hf: p1 = 12'd2372;
        endcase
    end

    always @ (*) begin
        case({ z_in[28], z_in[27], z_in[21], z_in[13] })
            4'h0: n0 = 12'd0;
            4'h1: n0 = 12'd990;
            4'h2: n0 = 12'd935;
            4'h3: n0 = 12'd1925;
            4'h4: n0 = 12'd157;
            4'h5: n0 = 12'd1147;
            4'h6: n0 = 12'd1092;
            4'h7: n0 = 12'd2082;
            4'h8: n0 = 12'd314;
            4'h9: n0 = 12'd1304;
            4'ha: n0 = 12'd1249;
            4'hb: n0 = 12'd2239;
            4'hc: n0 = 12'd471;
            4'hd: n0 = 12'd1461;
            4'he: n0 = 12'd1406;
            4'hf: n0 = 12'd2396;
        endcase
    end

    always @ (*) begin
        case({ z_in[31], z_in[24], z_in[20], z_in[19], z_in[16] })
            5'h00: n1 = 13'd0;
            5'h01: n1 = 13'd3329;
            5'h02: n1 = 13'd3677;
            5'h03: n1 = 13'd2415;
            5'h04: n1 = 13'd2763;
            5'h05: n1 = 13'd1501;
            5'h06: n1 = 13'd1849;
            5'h07: n1 = 13'd587;
            5'h08: n1 = 13'd2889;
            5'h09: n1 = 13'd1627;
            5'h0a: n1 = 13'd1975;
            5'h0b: n1 = 13'd713;
            5'h0c: n1 = 13'd1061;
            5'h0d: n1 = 13'd4390;
            5'h0e: n1 = 13'd147;
            5'h0f: n1 = 13'd3476;
            5'h10: n1 = 13'd2512;
            5'h11: n1 = 13'd1250;
            5'h12: n1 = 13'd1598;
            5'h13: n1 = 13'd336;
            5'h14: n1 = 13'd684;
            5'h15: n1 = 13'd4013;
            5'h16: n1 = 13'd4361;
            5'h17: n1 = 13'd3099;
            5'h18: n1 = 13'd810;
            5'h19: n1 = 13'd4139;
            5'h1a: n1 = 13'd4487;
            5'h1b: n1 = 13'd3225;
            5'h1c: n1 = 13'd3573;
            5'h1d: n1 = 13'd2311;
            5'h1e: n1 = 13'd2659;
            5'h1f: n1 = 13'd1397;
        endcase
    end

    always @ (*) begin
        case({ z_in[29], z_in[25], z_in[12] })
            3'h0: n2 = 12'd0;
            3'h1: n2 = 12'd495;
            3'h2: n2 = 12'd1187;
            3'h3: n2 = 12'd1682;
            3'h4: n2 = 12'd628;
            3'h5: n2 = 12'd1123;
            3'h6: n2 = 12'd1815;
            3'h7: n2 = 12'd2310;
        endcase
    end

    always @ (*) begin
        case({ z_in[30], z_in[26], z_in[22], z_in[17], z_in[14] })
            5'h00: n3 = 13'd0;
            5'h01: n3 = 13'd1980;
            5'h02: n3 = 13'd2067;
            5'h03: n3 = 13'd4047;
            5'h04: n3 = 13'd1870;
            5'h05: n3 = 13'd3850;
            5'h06: n3 = 13'd3937;
            5'h07: n3 = 13'd1326;
            5'h08: n3 = 13'd2374;
            5'h09: n3 = 13'd4354;
            5'h0a: n3 = 13'd4441;
            5'h0b: n3 = 13'd1830;
            5'h0c: n3 = 13'd4244;
            5'h0d: n3 = 13'd1633;
            5'h0e: n3 = 13'd1720;
            5'h0f: n3 = 13'd3700;
            5'h10: n3 = 13'd1256;
            5'h11: n3 = 13'd3236;
            5'h12: n3 = 13'd3323;
            5'h13: n3 = 13'd712;
            5'h14: n3 = 13'd3126;
            5'h15: n3 = 13'd515;
            5'h16: n3 = 13'd602;
            5'h17: n3 = 13'd2582;
            5'h18: n3 = 13'd3630;
            5'h19: n3 = 13'd1019;
            5'h1a: n3 = 13'd1106;
            5'h1b: n3 = 13'd3086;
            5'h1c: n3 = 13'd909;
            5'h1d: n3 = 13'd2889;
            5'h1e: n3 = 13'd2976;
            5'h1f: n3 = 13'd365;
        endcase
    end

endmodule
