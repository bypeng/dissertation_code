module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam B_LEN = 'd1815;
  localparam B_DEPTH = 'd11;
  localparam R_LEN = 'd1277;
  localparam R_DEPTH = 'd11;

  input              clk;
  input      [10: 0] in_addr;
  output reg [ 7: 0] in_data;
  input      [10: 0] out_addr;
  output reg [13: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      11'd0    : in_data <= 8'h08;
      11'd1    : in_data <= 8'h82;
      11'd2    : in_data <= 8'h6c;
      11'd3    : in_data <= 8'ha2;
      11'd4    : in_data <= 8'hc1;
      11'd5    : in_data <= 8'h89;
      11'd6    : in_data <= 8'hde;
      11'd7    : in_data <= 8'haa;
      11'd8    : in_data <= 8'h39;
      11'd9    : in_data <= 8'h2c;
      11'd10   : in_data <= 8'hc7;
      11'd11   : in_data <= 8'h6e;
      11'd12   : in_data <= 8'h21;
      11'd13   : in_data <= 8'h9b;
      11'd14   : in_data <= 8'hbe;
      11'd15   : in_data <= 8'h45;
      11'd16   : in_data <= 8'hbc;
      11'd17   : in_data <= 8'hb3;
      11'd18   : in_data <= 8'he9;
      11'd19   : in_data <= 8'heb;
      11'd20   : in_data <= 8'h49;
      11'd21   : in_data <= 8'hab;
      11'd22   : in_data <= 8'h06;
      11'd23   : in_data <= 8'h74;
      11'd24   : in_data <= 8'hf6;
      11'd25   : in_data <= 8'h5a;
      11'd26   : in_data <= 8'h75;
      11'd27   : in_data <= 8'hb4;
      11'd28   : in_data <= 8'h8e;
      11'd29   : in_data <= 8'hc2;
      11'd30   : in_data <= 8'hb2;
      11'd31   : in_data <= 8'h15;
      11'd32   : in_data <= 8'he5;
      11'd33   : in_data <= 8'h48;
      11'd34   : in_data <= 8'h36;
      11'd35   : in_data <= 8'h0b;
      11'd36   : in_data <= 8'h13;
      11'd37   : in_data <= 8'h03;
      11'd38   : in_data <= 8'h38;
      11'd39   : in_data <= 8'h56;
      11'd40   : in_data <= 8'ha0;
      11'd41   : in_data <= 8'hf3;
      11'd42   : in_data <= 8'hc9;
      11'd43   : in_data <= 8'h67;
      11'd44   : in_data <= 8'h86;
      11'd45   : in_data <= 8'hfa;
      11'd46   : in_data <= 8'h20;
      11'd47   : in_data <= 8'hd8;
      11'd48   : in_data <= 8'he5;
      11'd49   : in_data <= 8'haf;
      11'd50   : in_data <= 8'h87;
      11'd51   : in_data <= 8'h11;
      11'd52   : in_data <= 8'h35;
      11'd53   : in_data <= 8'h89;
      11'd54   : in_data <= 8'h90;
      11'd55   : in_data <= 8'h40;
      11'd56   : in_data <= 8'h70;
      11'd57   : in_data <= 8'h8e;
      11'd58   : in_data <= 8'h9a;
      11'd59   : in_data <= 8'h71;
      11'd60   : in_data <= 8'hd4;
      11'd61   : in_data <= 8'h2d;
      11'd62   : in_data <= 8'h74;
      11'd63   : in_data <= 8'h78;
      11'd64   : in_data <= 8'h50;
      11'd65   : in_data <= 8'h29;
      11'd66   : in_data <= 8'h38;
      11'd67   : in_data <= 8'h02;
      11'd68   : in_data <= 8'h4c;
      11'd69   : in_data <= 8'hee;
      11'd70   : in_data <= 8'h0b;
      11'd71   : in_data <= 8'h94;
      11'd72   : in_data <= 8'h26;
      11'd73   : in_data <= 8'h3e;
      11'd74   : in_data <= 8'h08;
      11'd75   : in_data <= 8'hc2;
      11'd76   : in_data <= 8'h45;
      11'd77   : in_data <= 8'h23;
      11'd78   : in_data <= 8'h88;
      11'd79   : in_data <= 8'hc6;
      11'd80   : in_data <= 8'hfa;
      11'd81   : in_data <= 8'h02;
      11'd82   : in_data <= 8'hda;
      11'd83   : in_data <= 8'h57;
      11'd84   : in_data <= 8'he0;
      11'd85   : in_data <= 8'hc7;
      11'd86   : in_data <= 8'h55;
      11'd87   : in_data <= 8'h5e;
      11'd88   : in_data <= 8'hc8;
      11'd89   : in_data <= 8'hcb;
      11'd90   : in_data <= 8'h71;
      11'd91   : in_data <= 8'h28;
      11'd92   : in_data <= 8'hf1;
      11'd93   : in_data <= 8'h67;
      11'd94   : in_data <= 8'hfb;
      11'd95   : in_data <= 8'h61;
      11'd96   : in_data <= 8'hd9;
      11'd97   : in_data <= 8'h8e;
      11'd98   : in_data <= 8'h35;
      11'd99   : in_data <= 8'h40;
      11'd100  : in_data <= 8'h5b;
      11'd101  : in_data <= 8'h78;
      11'd102  : in_data <= 8'h37;
      11'd103  : in_data <= 8'hf7;
      11'd104  : in_data <= 8'hbc;
      11'd105  : in_data <= 8'h10;
      11'd106  : in_data <= 8'hc3;
      11'd107  : in_data <= 8'h5e;
      11'd108  : in_data <= 8'hdc;
      11'd109  : in_data <= 8'h0c;
      11'd110  : in_data <= 8'hb3;
      11'd111  : in_data <= 8'h8c;
      11'd112  : in_data <= 8'h18;
      11'd113  : in_data <= 8'h82;
      11'd114  : in_data <= 8'h46;
      11'd115  : in_data <= 8'he5;
      11'd116  : in_data <= 8'h55;
      11'd117  : in_data <= 8'h51;
      11'd118  : in_data <= 8'h5d;
      11'd119  : in_data <= 8'hee;
      11'd120  : in_data <= 8'hbb;
      11'd121  : in_data <= 8'h6e;
      11'd122  : in_data <= 8'hf3;
      11'd123  : in_data <= 8'h9e;
      11'd124  : in_data <= 8'hb9;
      11'd125  : in_data <= 8'hed;
      11'd126  : in_data <= 8'hda;
      11'd127  : in_data <= 8'he9;
      11'd128  : in_data <= 8'h4a;
      11'd129  : in_data <= 8'h46;
      11'd130  : in_data <= 8'h46;
      11'd131  : in_data <= 8'h5b;
      11'd132  : in_data <= 8'h59;
      11'd133  : in_data <= 8'h0d;
      11'd134  : in_data <= 8'hd4;
      11'd135  : in_data <= 8'hea;
      11'd136  : in_data <= 8'hf9;
      11'd137  : in_data <= 8'h24;
      11'd138  : in_data <= 8'hb9;
      11'd139  : in_data <= 8'h03;
      11'd140  : in_data <= 8'h6f;
      11'd141  : in_data <= 8'h32;
      11'd142  : in_data <= 8'h90;
      11'd143  : in_data <= 8'h47;
      11'd144  : in_data <= 8'h83;
      11'd145  : in_data <= 8'h04;
      11'd146  : in_data <= 8'h77;
      11'd147  : in_data <= 8'heb;
      11'd148  : in_data <= 8'ha6;
      11'd149  : in_data <= 8'hf8;
      11'd150  : in_data <= 8'hb6;
      11'd151  : in_data <= 8'h6a;
      11'd152  : in_data <= 8'h75;
      11'd153  : in_data <= 8'h6f;
      11'd154  : in_data <= 8'he9;
      11'd155  : in_data <= 8'h62;
      11'd156  : in_data <= 8'hb8;
      11'd157  : in_data <= 8'hd4;
      11'd158  : in_data <= 8'hfa;
      11'd159  : in_data <= 8'hdd;
      11'd160  : in_data <= 8'hbc;
      11'd161  : in_data <= 8'hee;
      11'd162  : in_data <= 8'h0b;
      11'd163  : in_data <= 8'hdc;
      11'd164  : in_data <= 8'h8d;
      11'd165  : in_data <= 8'h11;
      11'd166  : in_data <= 8'h5f;
      11'd167  : in_data <= 8'h16;
      11'd168  : in_data <= 8'h64;
      11'd169  : in_data <= 8'hc2;
      11'd170  : in_data <= 8'ha1;
      11'd171  : in_data <= 8'h1f;
      11'd172  : in_data <= 8'hf2;
      11'd173  : in_data <= 8'hc8;
      11'd174  : in_data <= 8'h27;
      11'd175  : in_data <= 8'hd5;
      11'd176  : in_data <= 8'h21;
      11'd177  : in_data <= 8'hec;
      11'd178  : in_data <= 8'h2d;
      11'd179  : in_data <= 8'hfa;
      11'd180  : in_data <= 8'hef;
      11'd181  : in_data <= 8'hf2;
      11'd182  : in_data <= 8'h1d;
      11'd183  : in_data <= 8'hc8;
      11'd184  : in_data <= 8'he0;
      11'd185  : in_data <= 8'h71;
      11'd186  : in_data <= 8'hb6;
      11'd187  : in_data <= 8'he4;
      11'd188  : in_data <= 8'hce;
      11'd189  : in_data <= 8'h5e;
      11'd190  : in_data <= 8'h92;
      11'd191  : in_data <= 8'h29;
      11'd192  : in_data <= 8'ha9;
      11'd193  : in_data <= 8'h78;
      11'd194  : in_data <= 8'h29;
      11'd195  : in_data <= 8'h99;
      11'd196  : in_data <= 8'h55;
      11'd197  : in_data <= 8'h1f;
      11'd198  : in_data <= 8'h97;
      11'd199  : in_data <= 8'h4c;
      11'd200  : in_data <= 8'h3f;
      11'd201  : in_data <= 8'he3;
      11'd202  : in_data <= 8'h2e;
      11'd203  : in_data <= 8'ha1;
      11'd204  : in_data <= 8'h5c;
      11'd205  : in_data <= 8'h95;
      11'd206  : in_data <= 8'h29;
      11'd207  : in_data <= 8'h62;
      11'd208  : in_data <= 8'h1c;
      11'd209  : in_data <= 8'hdd;
      11'd210  : in_data <= 8'h5e;
      11'd211  : in_data <= 8'hfc;
      11'd212  : in_data <= 8'h36;
      11'd213  : in_data <= 8'h33;
      11'd214  : in_data <= 8'h64;
      11'd215  : in_data <= 8'hb3;
      11'd216  : in_data <= 8'h5e;
      11'd217  : in_data <= 8'h16;
      11'd218  : in_data <= 8'haa;
      11'd219  : in_data <= 8'h20;
      11'd220  : in_data <= 8'h93;
      11'd221  : in_data <= 8'hc7;
      11'd222  : in_data <= 8'h68;
      11'd223  : in_data <= 8'hda;
      11'd224  : in_data <= 8'h63;
      11'd225  : in_data <= 8'hc4;
      11'd226  : in_data <= 8'h24;
      11'd227  : in_data <= 8'h3a;
      11'd228  : in_data <= 8'h68;
      11'd229  : in_data <= 8'he3;
      11'd230  : in_data <= 8'hb3;
      11'd231  : in_data <= 8'h30;
      11'd232  : in_data <= 8'h07;
      11'd233  : in_data <= 8'he4;
      11'd234  : in_data <= 8'h97;
      11'd235  : in_data <= 8'h44;
      11'd236  : in_data <= 8'hdd;
      11'd237  : in_data <= 8'h88;
      11'd238  : in_data <= 8'he6;
      11'd239  : in_data <= 8'h84;
      11'd240  : in_data <= 8'h1c;
      11'd241  : in_data <= 8'h55;
      11'd242  : in_data <= 8'hb8;
      11'd243  : in_data <= 8'h32;
      11'd244  : in_data <= 8'hcb;
      11'd245  : in_data <= 8'hdc;
      11'd246  : in_data <= 8'hb3;
      11'd247  : in_data <= 8'h50;
      11'd248  : in_data <= 8'h63;
      11'd249  : in_data <= 8'hf2;
      11'd250  : in_data <= 8'hda;
      11'd251  : in_data <= 8'h87;
      11'd252  : in_data <= 8'hf9;
      11'd253  : in_data <= 8'h06;
      11'd254  : in_data <= 8'h4b;
      11'd255  : in_data <= 8'h3f;
      11'd256  : in_data <= 8'h2f;
      11'd257  : in_data <= 8'hd1;
      11'd258  : in_data <= 8'h4a;
      11'd259  : in_data <= 8'hf2;
      11'd260  : in_data <= 8'hec;
      11'd261  : in_data <= 8'h4a;
      11'd262  : in_data <= 8'h98;
      11'd263  : in_data <= 8'hc0;
      11'd264  : in_data <= 8'h06;
      11'd265  : in_data <= 8'h24;
      11'd266  : in_data <= 8'h25;
      11'd267  : in_data <= 8'h12;
      11'd268  : in_data <= 8'h82;
      11'd269  : in_data <= 8'h09;
      11'd270  : in_data <= 8'h40;
      11'd271  : in_data <= 8'hcb;
      11'd272  : in_data <= 8'h9f;
      11'd273  : in_data <= 8'h5d;
      11'd274  : in_data <= 8'h47;
      11'd275  : in_data <= 8'h77;
      11'd276  : in_data <= 8'h02;
      11'd277  : in_data <= 8'h30;
      11'd278  : in_data <= 8'h8d;
      11'd279  : in_data <= 8'hf1;
      11'd280  : in_data <= 8'h19;
      11'd281  : in_data <= 8'hd6;
      11'd282  : in_data <= 8'ha6;
      11'd283  : in_data <= 8'h15;
      11'd284  : in_data <= 8'ha5;
      11'd285  : in_data <= 8'hc9;
      11'd286  : in_data <= 8'h93;
      11'd287  : in_data <= 8'h3c;
      11'd288  : in_data <= 8'hca;
      11'd289  : in_data <= 8'h89;
      11'd290  : in_data <= 8'h15;
      11'd291  : in_data <= 8'h9b;
      11'd292  : in_data <= 8'h34;
      11'd293  : in_data <= 8'hb8;
      11'd294  : in_data <= 8'hb7;
      11'd295  : in_data <= 8'h36;
      11'd296  : in_data <= 8'h5d;
      11'd297  : in_data <= 8'h3d;
      11'd298  : in_data <= 8'h30;
      11'd299  : in_data <= 8'h4e;
      11'd300  : in_data <= 8'h53;
      11'd301  : in_data <= 8'h63;
      11'd302  : in_data <= 8'h02;
      11'd303  : in_data <= 8'h97;
      11'd304  : in_data <= 8'h12;
      11'd305  : in_data <= 8'h5b;
      11'd306  : in_data <= 8'h17;
      11'd307  : in_data <= 8'h8e;
      11'd308  : in_data <= 8'hf0;
      11'd309  : in_data <= 8'h2f;
      11'd310  : in_data <= 8'h37;
      11'd311  : in_data <= 8'h9b;
      11'd312  : in_data <= 8'h48;
      11'd313  : in_data <= 8'h2a;
      11'd314  : in_data <= 8'h8d;
      11'd315  : in_data <= 8'he9;
      11'd316  : in_data <= 8'h4a;
      11'd317  : in_data <= 8'h83;
      11'd318  : in_data <= 8'hc1;
      11'd319  : in_data <= 8'h63;
      11'd320  : in_data <= 8'h8d;
      11'd321  : in_data <= 8'h47;
      11'd322  : in_data <= 8'h15;
      11'd323  : in_data <= 8'h94;
      11'd324  : in_data <= 8'hf1;
      11'd325  : in_data <= 8'hc9;
      11'd326  : in_data <= 8'h20;
      11'd327  : in_data <= 8'h01;
      11'd328  : in_data <= 8'h39;
      11'd329  : in_data <= 8'hab;
      11'd330  : in_data <= 8'h55;
      11'd331  : in_data <= 8'hdc;
      11'd332  : in_data <= 8'h12;
      11'd333  : in_data <= 8'h91;
      11'd334  : in_data <= 8'h68;
      11'd335  : in_data <= 8'h20;
      11'd336  : in_data <= 8'h6c;
      11'd337  : in_data <= 8'h35;
      11'd338  : in_data <= 8'h9f;
      11'd339  : in_data <= 8'he6;
      11'd340  : in_data <= 8'h51;
      11'd341  : in_data <= 8'h60;
      11'd342  : in_data <= 8'hc2;
      11'd343  : in_data <= 8'hc7;
      11'd344  : in_data <= 8'h19;
      11'd345  : in_data <= 8'hf4;
      11'd346  : in_data <= 8'h5e;
      11'd347  : in_data <= 8'h1c;
      11'd348  : in_data <= 8'h46;
      11'd349  : in_data <= 8'h73;
      11'd350  : in_data <= 8'h2c;
      11'd351  : in_data <= 8'h50;
      11'd352  : in_data <= 8'hcc;
      11'd353  : in_data <= 8'haf;
      11'd354  : in_data <= 8'hb8;
      11'd355  : in_data <= 8'hc3;
      11'd356  : in_data <= 8'h2f;
      11'd357  : in_data <= 8'h6d;
      11'd358  : in_data <= 8'h12;
      11'd359  : in_data <= 8'hd0;
      11'd360  : in_data <= 8'ha9;
      11'd361  : in_data <= 8'hbf;
      11'd362  : in_data <= 8'h36;
      11'd363  : in_data <= 8'hd7;
      11'd364  : in_data <= 8'h5e;
      11'd365  : in_data <= 8'h0c;
      11'd366  : in_data <= 8'h39;
      11'd367  : in_data <= 8'h3b;
      11'd368  : in_data <= 8'h4f;
      11'd369  : in_data <= 8'h35;
      11'd370  : in_data <= 8'h51;
      11'd371  : in_data <= 8'h16;
      11'd372  : in_data <= 8'hb4;
      11'd373  : in_data <= 8'h76;
      11'd374  : in_data <= 8'h49;
      11'd375  : in_data <= 8'h23;
      11'd376  : in_data <= 8'h15;
      11'd377  : in_data <= 8'h27;
      11'd378  : in_data <= 8'h73;
      11'd379  : in_data <= 8'hba;
      11'd380  : in_data <= 8'h84;
      11'd381  : in_data <= 8'he3;
      11'd382  : in_data <= 8'h58;
      11'd383  : in_data <= 8'hef;
      11'd384  : in_data <= 8'hdb;
      11'd385  : in_data <= 8'h83;
      11'd386  : in_data <= 8'hd0;
      11'd387  : in_data <= 8'h56;
      11'd388  : in_data <= 8'h83;
      11'd389  : in_data <= 8'h72;
      11'd390  : in_data <= 8'h4f;
      11'd391  : in_data <= 8'hcf;
      11'd392  : in_data <= 8'hf1;
      11'd393  : in_data <= 8'h03;
      11'd394  : in_data <= 8'hfb;
      11'd395  : in_data <= 8'he5;
      11'd396  : in_data <= 8'heb;
      11'd397  : in_data <= 8'h70;
      11'd398  : in_data <= 8'hcb;
      11'd399  : in_data <= 8'hb6;
      11'd400  : in_data <= 8'hfc;
      11'd401  : in_data <= 8'h26;
      11'd402  : in_data <= 8'h62;
      11'd403  : in_data <= 8'h7c;
      11'd404  : in_data <= 8'h05;
      11'd405  : in_data <= 8'h3a;
      11'd406  : in_data <= 8'h79;
      11'd407  : in_data <= 8'h7d;
      11'd408  : in_data <= 8'hc8;
      11'd409  : in_data <= 8'h11;
      11'd410  : in_data <= 8'h6e;
      11'd411  : in_data <= 8'hda;
      11'd412  : in_data <= 8'h25;
      11'd413  : in_data <= 8'h1a;
      11'd414  : in_data <= 8'h35;
      11'd415  : in_data <= 8'h23;
      11'd416  : in_data <= 8'h4c;
      11'd417  : in_data <= 8'h84;
      11'd418  : in_data <= 8'h89;
      11'd419  : in_data <= 8'hb4;
      11'd420  : in_data <= 8'he0;
      11'd421  : in_data <= 8'h7f;
      11'd422  : in_data <= 8'h60;
      11'd423  : in_data <= 8'h9a;
      11'd424  : in_data <= 8'h84;
      11'd425  : in_data <= 8'hf2;
      11'd426  : in_data <= 8'h57;
      11'd427  : in_data <= 8'hb9;
      11'd428  : in_data <= 8'h1f;
      11'd429  : in_data <= 8'h39;
      11'd430  : in_data <= 8'hec;
      11'd431  : in_data <= 8'h4d;
      11'd432  : in_data <= 8'he3;
      11'd433  : in_data <= 8'h61;
      11'd434  : in_data <= 8'hc1;
      11'd435  : in_data <= 8'h2f;
      11'd436  : in_data <= 8'hbb;
      11'd437  : in_data <= 8'h08;
      11'd438  : in_data <= 8'hd3;
      11'd439  : in_data <= 8'h0c;
      11'd440  : in_data <= 8'h3e;
      11'd441  : in_data <= 8'hf7;
      11'd442  : in_data <= 8'h18;
      11'd443  : in_data <= 8'hf8;
      11'd444  : in_data <= 8'h62;
      11'd445  : in_data <= 8'ha0;
      11'd446  : in_data <= 8'h30;
      11'd447  : in_data <= 8'h4f;
      11'd448  : in_data <= 8'h4e;
      11'd449  : in_data <= 8'hb7;
      11'd450  : in_data <= 8'h84;
      11'd451  : in_data <= 8'h24;
      11'd452  : in_data <= 8'hc7;
      11'd453  : in_data <= 8'hae;
      11'd454  : in_data <= 8'h2c;
      11'd455  : in_data <= 8'hc1;
      11'd456  : in_data <= 8'hcc;
      11'd457  : in_data <= 8'h38;
      11'd458  : in_data <= 8'h67;
      11'd459  : in_data <= 8'h5e;
      11'd460  : in_data <= 8'h88;
      11'd461  : in_data <= 8'h2b;
      11'd462  : in_data <= 8'hac;
      11'd463  : in_data <= 8'he9;
      11'd464  : in_data <= 8'hcc;
      11'd465  : in_data <= 8'h45;
      11'd466  : in_data <= 8'h59;
      11'd467  : in_data <= 8'h45;
      11'd468  : in_data <= 8'hbc;
      11'd469  : in_data <= 8'h3a;
      11'd470  : in_data <= 8'h43;
      11'd471  : in_data <= 8'h75;
      11'd472  : in_data <= 8'h83;
      11'd473  : in_data <= 8'h74;
      11'd474  : in_data <= 8'h09;
      11'd475  : in_data <= 8'h80;
      11'd476  : in_data <= 8'h7b;
      11'd477  : in_data <= 8'h2b;
      11'd478  : in_data <= 8'h6e;
      11'd479  : in_data <= 8'h43;
      11'd480  : in_data <= 8'h2d;
      11'd481  : in_data <= 8'h9c;
      11'd482  : in_data <= 8'h85;
      11'd483  : in_data <= 8'hf1;
      11'd484  : in_data <= 8'he2;
      11'd485  : in_data <= 8'h22;
      11'd486  : in_data <= 8'h30;
      11'd487  : in_data <= 8'hd9;
      11'd488  : in_data <= 8'hd7;
      11'd489  : in_data <= 8'hed;
      11'd490  : in_data <= 8'hc0;
      11'd491  : in_data <= 8'hc6;
      11'd492  : in_data <= 8'he4;
      11'd493  : in_data <= 8'h5f;
      11'd494  : in_data <= 8'h24;
      11'd495  : in_data <= 8'h5f;
      11'd496  : in_data <= 8'hc0;
      11'd497  : in_data <= 8'hd7;
      11'd498  : in_data <= 8'hc9;
      11'd499  : in_data <= 8'h93;
      11'd500  : in_data <= 8'h6e;
      11'd501  : in_data <= 8'h00;
      11'd502  : in_data <= 8'hc2;
      11'd503  : in_data <= 8'h6c;
      11'd504  : in_data <= 8'h27;
      11'd505  : in_data <= 8'hb4;
      11'd506  : in_data <= 8'h65;
      11'd507  : in_data <= 8'had;
      11'd508  : in_data <= 8'h97;
      11'd509  : in_data <= 8'h79;
      11'd510  : in_data <= 8'hac;
      11'd511  : in_data <= 8'h51;
      11'd512  : in_data <= 8'hef;
      11'd513  : in_data <= 8'h11;
      11'd514  : in_data <= 8'ha1;
      11'd515  : in_data <= 8'h83;
      11'd516  : in_data <= 8'h3b;
      11'd517  : in_data <= 8'hd7;
      11'd518  : in_data <= 8'hb3;
      11'd519  : in_data <= 8'h5c;
      11'd520  : in_data <= 8'ha9;
      11'd521  : in_data <= 8'h80;
      11'd522  : in_data <= 8'hf8;
      11'd523  : in_data <= 8'h05;
      11'd524  : in_data <= 8'hec;
      11'd525  : in_data <= 8'hc8;
      11'd526  : in_data <= 8'hd5;
      11'd527  : in_data <= 8'h18;
      11'd528  : in_data <= 8'h6c;
      11'd529  : in_data <= 8'hfc;
      11'd530  : in_data <= 8'h8b;
      11'd531  : in_data <= 8'h3f;
      11'd532  : in_data <= 8'ha7;
      11'd533  : in_data <= 8'h7d;
      11'd534  : in_data <= 8'ha2;
      11'd535  : in_data <= 8'h42;
      11'd536  : in_data <= 8'h07;
      11'd537  : in_data <= 8'hec;
      11'd538  : in_data <= 8'ha9;
      11'd539  : in_data <= 8'h33;
      11'd540  : in_data <= 8'hf9;
      11'd541  : in_data <= 8'h7e;
      11'd542  : in_data <= 8'h8b;
      11'd543  : in_data <= 8'hb2;
      11'd544  : in_data <= 8'h9b;
      11'd545  : in_data <= 8'hd8;
      11'd546  : in_data <= 8'hae;
      11'd547  : in_data <= 8'haf;
      11'd548  : in_data <= 8'h92;
      11'd549  : in_data <= 8'ha7;
      11'd550  : in_data <= 8'hc7;
      11'd551  : in_data <= 8'h53;
      11'd552  : in_data <= 8'h45;
      11'd553  : in_data <= 8'h8f;
      11'd554  : in_data <= 8'hc1;
      11'd555  : in_data <= 8'h6b;
      11'd556  : in_data <= 8'he9;
      11'd557  : in_data <= 8'hb8;
      11'd558  : in_data <= 8'h13;
      11'd559  : in_data <= 8'h1b;
      11'd560  : in_data <= 8'hcf;
      11'd561  : in_data <= 8'hfd;
      11'd562  : in_data <= 8'h73;
      11'd563  : in_data <= 8'ha8;
      11'd564  : in_data <= 8'h59;
      11'd565  : in_data <= 8'hdd;
      11'd566  : in_data <= 8'hfc;
      11'd567  : in_data <= 8'h51;
      11'd568  : in_data <= 8'h02;
      11'd569  : in_data <= 8'hf8;
      11'd570  : in_data <= 8'h09;
      11'd571  : in_data <= 8'hf3;
      11'd572  : in_data <= 8'heb;
      11'd573  : in_data <= 8'he1;
      11'd574  : in_data <= 8'h93;
      11'd575  : in_data <= 8'hfb;
      11'd576  : in_data <= 8'hd5;
      11'd577  : in_data <= 8'h80;
      11'd578  : in_data <= 8'hde;
      11'd579  : in_data <= 8'he6;
      11'd580  : in_data <= 8'hf9;
      11'd581  : in_data <= 8'h0b;
      11'd582  : in_data <= 8'hdb;
      11'd583  : in_data <= 8'h5a;
      11'd584  : in_data <= 8'h36;
      11'd585  : in_data <= 8'hbb;
      11'd586  : in_data <= 8'h43;
      11'd587  : in_data <= 8'hf2;
      11'd588  : in_data <= 8'h64;
      11'd589  : in_data <= 8'h62;
      11'd590  : in_data <= 8'ha5;
      11'd591  : in_data <= 8'hc8;
      11'd592  : in_data <= 8'h55;
      11'd593  : in_data <= 8'h7f;
      11'd594  : in_data <= 8'h18;
      11'd595  : in_data <= 8'hdb;
      11'd596  : in_data <= 8'h75;
      11'd597  : in_data <= 8'hcf;
      11'd598  : in_data <= 8'h8a;
      11'd599  : in_data <= 8'h6b;
      11'd600  : in_data <= 8'h15;
      11'd601  : in_data <= 8'h85;
      11'd602  : in_data <= 8'h9d;
      11'd603  : in_data <= 8'h08;
      11'd604  : in_data <= 8'h55;
      11'd605  : in_data <= 8'hd8;
      11'd606  : in_data <= 8'h18;
      11'd607  : in_data <= 8'h50;
      11'd608  : in_data <= 8'h99;
      11'd609  : in_data <= 8'h88;
      11'd610  : in_data <= 8'hc9;
      11'd611  : in_data <= 8'h37;
      11'd612  : in_data <= 8'h64;
      11'd613  : in_data <= 8'hb6;
      11'd614  : in_data <= 8'h55;
      11'd615  : in_data <= 8'hb5;
      11'd616  : in_data <= 8'h6b;
      11'd617  : in_data <= 8'h03;
      11'd618  : in_data <= 8'h02;
      11'd619  : in_data <= 8'h32;
      11'd620  : in_data <= 8'h49;
      11'd621  : in_data <= 8'hfc;
      11'd622  : in_data <= 8'hdb;
      11'd623  : in_data <= 8'h7d;
      11'd624  : in_data <= 8'h00;
      11'd625  : in_data <= 8'h36;
      11'd626  : in_data <= 8'h94;
      11'd627  : in_data <= 8'hd6;
      11'd628  : in_data <= 8'h71;
      11'd629  : in_data <= 8'h16;
      11'd630  : in_data <= 8'h9b;
      11'd631  : in_data <= 8'h68;
      11'd632  : in_data <= 8'h51;
      11'd633  : in_data <= 8'he4;
      11'd634  : in_data <= 8'h48;
      11'd635  : in_data <= 8'h19;
      11'd636  : in_data <= 8'had;
      11'd637  : in_data <= 8'h6d;
      11'd638  : in_data <= 8'hd7;
      11'd639  : in_data <= 8'h86;
      11'd640  : in_data <= 8'hbe;
      11'd641  : in_data <= 8'hbb;
      11'd642  : in_data <= 8'hff;
      11'd643  : in_data <= 8'h98;
      11'd644  : in_data <= 8'hf3;
      11'd645  : in_data <= 8'h2b;
      11'd646  : in_data <= 8'h0c;
      11'd647  : in_data <= 8'he0;
      11'd648  : in_data <= 8'hec;
      11'd649  : in_data <= 8'hec;
      11'd650  : in_data <= 8'h26;
      11'd651  : in_data <= 8'h99;
      11'd652  : in_data <= 8'h53;
      11'd653  : in_data <= 8'h45;
      11'd654  : in_data <= 8'h98;
      11'd655  : in_data <= 8'h7b;
      11'd656  : in_data <= 8'h7e;
      11'd657  : in_data <= 8'h1e;
      11'd658  : in_data <= 8'hc9;
      11'd659  : in_data <= 8'hea;
      11'd660  : in_data <= 8'h9f;
      11'd661  : in_data <= 8'h0e;
      11'd662  : in_data <= 8'h8b;
      11'd663  : in_data <= 8'h88;
      11'd664  : in_data <= 8'h4f;
      11'd665  : in_data <= 8'h48;
      11'd666  : in_data <= 8'h58;
      11'd667  : in_data <= 8'h4d;
      11'd668  : in_data <= 8'h0c;
      11'd669  : in_data <= 8'hed;
      11'd670  : in_data <= 8'h43;
      11'd671  : in_data <= 8'h77;
      11'd672  : in_data <= 8'h75;
      11'd673  : in_data <= 8'h12;
      11'd674  : in_data <= 8'h1d;
      11'd675  : in_data <= 8'h04;
      11'd676  : in_data <= 8'hce;
      11'd677  : in_data <= 8'hbc;
      11'd678  : in_data <= 8'h50;
      11'd679  : in_data <= 8'h2b;
      11'd680  : in_data <= 8'h5b;
      11'd681  : in_data <= 8'h3d;
      11'd682  : in_data <= 8'hb8;
      11'd683  : in_data <= 8'h19;
      11'd684  : in_data <= 8'h07;
      11'd685  : in_data <= 8'ha0;
      11'd686  : in_data <= 8'h1e;
      11'd687  : in_data <= 8'h97;
      11'd688  : in_data <= 8'hd1;
      11'd689  : in_data <= 8'h28;
      11'd690  : in_data <= 8'h02;
      11'd691  : in_data <= 8'h24;
      11'd692  : in_data <= 8'h79;
      11'd693  : in_data <= 8'h52;
      11'd694  : in_data <= 8'he2;
      11'd695  : in_data <= 8'h10;
      11'd696  : in_data <= 8'hf5;
      11'd697  : in_data <= 8'hc2;
      11'd698  : in_data <= 8'h61;
      11'd699  : in_data <= 8'h10;
      11'd700  : in_data <= 8'hcf;
      11'd701  : in_data <= 8'h8d;
      11'd702  : in_data <= 8'h29;
      11'd703  : in_data <= 8'h5d;
      11'd704  : in_data <= 8'he4;
      11'd705  : in_data <= 8'he1;
      11'd706  : in_data <= 8'h6b;
      11'd707  : in_data <= 8'h4c;
      11'd708  : in_data <= 8'hf5;
      11'd709  : in_data <= 8'h49;
      11'd710  : in_data <= 8'hf4;
      11'd711  : in_data <= 8'h2e;
      11'd712  : in_data <= 8'h8e;
      11'd713  : in_data <= 8'he0;
      11'd714  : in_data <= 8'h1f;
      11'd715  : in_data <= 8'h8a;
      11'd716  : in_data <= 8'hce;
      11'd717  : in_data <= 8'h72;
      11'd718  : in_data <= 8'hfd;
      11'd719  : in_data <= 8'hfd;
      11'd720  : in_data <= 8'hdc;
      11'd721  : in_data <= 8'hf9;
      11'd722  : in_data <= 8'hc8;
      11'd723  : in_data <= 8'hec;
      11'd724  : in_data <= 8'hc0;
      11'd725  : in_data <= 8'hea;
      11'd726  : in_data <= 8'h04;
      11'd727  : in_data <= 8'ha3;
      11'd728  : in_data <= 8'hbd;
      11'd729  : in_data <= 8'h66;
      11'd730  : in_data <= 8'h95;
      11'd731  : in_data <= 8'h71;
      11'd732  : in_data <= 8'hf6;
      11'd733  : in_data <= 8'h6d;
      11'd734  : in_data <= 8'he1;
      11'd735  : in_data <= 8'h0e;
      11'd736  : in_data <= 8'h2e;
      11'd737  : in_data <= 8'h79;
      11'd738  : in_data <= 8'h3b;
      11'd739  : in_data <= 8'he0;
      11'd740  : in_data <= 8'haf;
      11'd741  : in_data <= 8'hcf;
      11'd742  : in_data <= 8'h24;
      11'd743  : in_data <= 8'h60;
      11'd744  : in_data <= 8'h7d;
      11'd745  : in_data <= 8'hc2;
      11'd746  : in_data <= 8'h90;
      11'd747  : in_data <= 8'hd5;
      11'd748  : in_data <= 8'h79;
      11'd749  : in_data <= 8'h91;
      11'd750  : in_data <= 8'hc5;
      11'd751  : in_data <= 8'h22;
      11'd752  : in_data <= 8'h2c;
      11'd753  : in_data <= 8'h91;
      11'd754  : in_data <= 8'hed;
      11'd755  : in_data <= 8'h12;
      11'd756  : in_data <= 8'h21;
      11'd757  : in_data <= 8'h81;
      11'd758  : in_data <= 8'h6d;
      11'd759  : in_data <= 8'h2e;
      11'd760  : in_data <= 8'hc2;
      11'd761  : in_data <= 8'he4;
      11'd762  : in_data <= 8'hcc;
      11'd763  : in_data <= 8'h63;
      11'd764  : in_data <= 8'h6c;
      11'd765  : in_data <= 8'h40;
      11'd766  : in_data <= 8'h23;
      11'd767  : in_data <= 8'hca;
      11'd768  : in_data <= 8'h8b;
      11'd769  : in_data <= 8'h5a;
      11'd770  : in_data <= 8'he0;
      11'd771  : in_data <= 8'h7c;
      11'd772  : in_data <= 8'h10;
      11'd773  : in_data <= 8'haa;
      11'd774  : in_data <= 8'h1e;
      11'd775  : in_data <= 8'h26;
      11'd776  : in_data <= 8'h1e;
      11'd777  : in_data <= 8'h8e;
      11'd778  : in_data <= 8'h41;
      11'd779  : in_data <= 8'hc2;
      11'd780  : in_data <= 8'h55;
      11'd781  : in_data <= 8'hbe;
      11'd782  : in_data <= 8'he5;
      11'd783  : in_data <= 8'ha0;
      11'd784  : in_data <= 8'h56;
      11'd785  : in_data <= 8'hd0;
      11'd786  : in_data <= 8'h65;
      11'd787  : in_data <= 8'h9a;
      11'd788  : in_data <= 8'hac;
      11'd789  : in_data <= 8'h8a;
      11'd790  : in_data <= 8'hb6;
      11'd791  : in_data <= 8'h06;
      11'd792  : in_data <= 8'hea;
      11'd793  : in_data <= 8'hd0;
      11'd794  : in_data <= 8'h43;
      11'd795  : in_data <= 8'h2e;
      11'd796  : in_data <= 8'hff;
      11'd797  : in_data <= 8'h0b;
      11'd798  : in_data <= 8'hdb;
      11'd799  : in_data <= 8'h54;
      11'd800  : in_data <= 8'h54;
      11'd801  : in_data <= 8'h7b;
      11'd802  : in_data <= 8'hc3;
      11'd803  : in_data <= 8'hc2;
      11'd804  : in_data <= 8'hbb;
      11'd805  : in_data <= 8'h90;
      11'd806  : in_data <= 8'he8;
      11'd807  : in_data <= 8'hd6;
      11'd808  : in_data <= 8'hf5;
      11'd809  : in_data <= 8'h9f;
      11'd810  : in_data <= 8'hb4;
      11'd811  : in_data <= 8'h20;
      11'd812  : in_data <= 8'hd4;
      11'd813  : in_data <= 8'h4f;
      11'd814  : in_data <= 8'h16;
      11'd815  : in_data <= 8'h3d;
      11'd816  : in_data <= 8'hfe;
      11'd817  : in_data <= 8'h6e;
      11'd818  : in_data <= 8'h40;
      11'd819  : in_data <= 8'h65;
      11'd820  : in_data <= 8'h59;
      11'd821  : in_data <= 8'h95;
      11'd822  : in_data <= 8'he7;
      11'd823  : in_data <= 8'h30;
      11'd824  : in_data <= 8'h11;
      11'd825  : in_data <= 8'haf;
      11'd826  : in_data <= 8'hd7;
      11'd827  : in_data <= 8'hff;
      11'd828  : in_data <= 8'ha3;
      11'd829  : in_data <= 8'h43;
      11'd830  : in_data <= 8'h1f;
      11'd831  : in_data <= 8'hf5;
      11'd832  : in_data <= 8'h69;
      11'd833  : in_data <= 8'hbb;
      11'd834  : in_data <= 8'h33;
      11'd835  : in_data <= 8'hf8;
      11'd836  : in_data <= 8'hc5;
      11'd837  : in_data <= 8'h28;
      11'd838  : in_data <= 8'haf;
      11'd839  : in_data <= 8'h76;
      11'd840  : in_data <= 8'he3;
      11'd841  : in_data <= 8'h8e;
      11'd842  : in_data <= 8'h25;
      11'd843  : in_data <= 8'he1;
      11'd844  : in_data <= 8'h53;
      11'd845  : in_data <= 8'hd7;
      11'd846  : in_data <= 8'hf5;
      11'd847  : in_data <= 8'h67;
      11'd848  : in_data <= 8'h6b;
      11'd849  : in_data <= 8'h41;
      11'd850  : in_data <= 8'h5d;
      11'd851  : in_data <= 8'hc9;
      11'd852  : in_data <= 8'h02;
      11'd853  : in_data <= 8'h7a;
      11'd854  : in_data <= 8'h9e;
      11'd855  : in_data <= 8'hb0;
      11'd856  : in_data <= 8'h43;
      11'd857  : in_data <= 8'hd7;
      11'd858  : in_data <= 8'h2f;
      11'd859  : in_data <= 8'ha3;
      11'd860  : in_data <= 8'h13;
      11'd861  : in_data <= 8'h07;
      11'd862  : in_data <= 8'h25;
      11'd863  : in_data <= 8'hd9;
      11'd864  : in_data <= 8'h67;
      11'd865  : in_data <= 8'haa;
      11'd866  : in_data <= 8'hee;
      11'd867  : in_data <= 8'h64;
      11'd868  : in_data <= 8'h67;
      11'd869  : in_data <= 8'ha0;
      11'd870  : in_data <= 8'h29;
      11'd871  : in_data <= 8'he3;
      11'd872  : in_data <= 8'hb1;
      11'd873  : in_data <= 8'h6b;
      11'd874  : in_data <= 8'hd8;
      11'd875  : in_data <= 8'he7;
      11'd876  : in_data <= 8'h41;
      11'd877  : in_data <= 8'h2f;
      11'd878  : in_data <= 8'h2d;
      11'd879  : in_data <= 8'he2;
      11'd880  : in_data <= 8'h68;
      11'd881  : in_data <= 8'hcc;
      11'd882  : in_data <= 8'hcf;
      11'd883  : in_data <= 8'hf2;
      11'd884  : in_data <= 8'hf3;
      11'd885  : in_data <= 8'h45;
      11'd886  : in_data <= 8'h3b;
      11'd887  : in_data <= 8'h22;
      11'd888  : in_data <= 8'he3;
      11'd889  : in_data <= 8'h36;
      11'd890  : in_data <= 8'hb1;
      11'd891  : in_data <= 8'h50;
      11'd892  : in_data <= 8'h16;
      11'd893  : in_data <= 8'h75;
      11'd894  : in_data <= 8'hf8;
      11'd895  : in_data <= 8'h40;
      11'd896  : in_data <= 8'hec;
      11'd897  : in_data <= 8'had;
      11'd898  : in_data <= 8'h13;
      11'd899  : in_data <= 8'hf5;
      11'd900  : in_data <= 8'h66;
      11'd901  : in_data <= 8'h73;
      11'd902  : in_data <= 8'hc5;
      11'd903  : in_data <= 8'h75;
      11'd904  : in_data <= 8'h50;
      11'd905  : in_data <= 8'h5b;
      11'd906  : in_data <= 8'hd1;
      11'd907  : in_data <= 8'h59;
      11'd908  : in_data <= 8'h92;
      11'd909  : in_data <= 8'ha0;
      11'd910  : in_data <= 8'hef;
      11'd911  : in_data <= 8'he6;
      11'd912  : in_data <= 8'h4c;
      11'd913  : in_data <= 8'h90;
      11'd914  : in_data <= 8'hd8;
      11'd915  : in_data <= 8'hb4;
      11'd916  : in_data <= 8'h14;
      11'd917  : in_data <= 8'h38;
      11'd918  : in_data <= 8'h23;
      11'd919  : in_data <= 8'ha3;
      11'd920  : in_data <= 8'h42;
      11'd921  : in_data <= 8'hfe;
      11'd922  : in_data <= 8'hef;
      11'd923  : in_data <= 8'ha3;
      11'd924  : in_data <= 8'h5a;
      11'd925  : in_data <= 8'h12;
      11'd926  : in_data <= 8'hb6;
      11'd927  : in_data <= 8'h9b;
      11'd928  : in_data <= 8'h30;
      11'd929  : in_data <= 8'h25;
      11'd930  : in_data <= 8'h5a;
      11'd931  : in_data <= 8'h5d;
      11'd932  : in_data <= 8'hff;
      11'd933  : in_data <= 8'hee;
      11'd934  : in_data <= 8'h4c;
      11'd935  : in_data <= 8'h1d;
      11'd936  : in_data <= 8'h2b;
      11'd937  : in_data <= 8'h35;
      11'd938  : in_data <= 8'h71;
      11'd939  : in_data <= 8'ha7;
      11'd940  : in_data <= 8'he7;
      11'd941  : in_data <= 8'h33;
      11'd942  : in_data <= 8'hcd;
      11'd943  : in_data <= 8'h25;
      11'd944  : in_data <= 8'h17;
      11'd945  : in_data <= 8'had;
      11'd946  : in_data <= 8'hf1;
      11'd947  : in_data <= 8'he0;
      11'd948  : in_data <= 8'h39;
      11'd949  : in_data <= 8'h3a;
      11'd950  : in_data <= 8'h27;
      11'd951  : in_data <= 8'h73;
      11'd952  : in_data <= 8'hc9;
      11'd953  : in_data <= 8'h09;
      11'd954  : in_data <= 8'h91;
      11'd955  : in_data <= 8'hab;
      11'd956  : in_data <= 8'hf7;
      11'd957  : in_data <= 8'h02;
      11'd958  : in_data <= 8'h81;
      11'd959  : in_data <= 8'h75;
      11'd960  : in_data <= 8'h93;
      11'd961  : in_data <= 8'h46;
      11'd962  : in_data <= 8'hf3;
      11'd963  : in_data <= 8'hc7;
      11'd964  : in_data <= 8'h74;
      11'd965  : in_data <= 8'h81;
      11'd966  : in_data <= 8'h08;
      11'd967  : in_data <= 8'hc9;
      11'd968  : in_data <= 8'h61;
      11'd969  : in_data <= 8'h47;
      11'd970  : in_data <= 8'hca;
      11'd971  : in_data <= 8'h01;
      11'd972  : in_data <= 8'h92;
      11'd973  : in_data <= 8'hcb;
      11'd974  : in_data <= 8'h14;
      11'd975  : in_data <= 8'hb1;
      11'd976  : in_data <= 8'hea;
      11'd977  : in_data <= 8'h03;
      11'd978  : in_data <= 8'h1a;
      11'd979  : in_data <= 8'hb1;
      11'd980  : in_data <= 8'hdd;
      11'd981  : in_data <= 8'h4f;
      11'd982  : in_data <= 8'h26;
      11'd983  : in_data <= 8'h57;
      11'd984  : in_data <= 8'h42;
      11'd985  : in_data <= 8'he8;
      11'd986  : in_data <= 8'ha3;
      11'd987  : in_data <= 8'h20;
      11'd988  : in_data <= 8'hd5;
      11'd989  : in_data <= 8'h2a;
      11'd990  : in_data <= 8'h06;
      11'd991  : in_data <= 8'h15;
      11'd992  : in_data <= 8'h53;
      11'd993  : in_data <= 8'h0e;
      11'd994  : in_data <= 8'hf0;
      11'd995  : in_data <= 8'h5a;
      11'd996  : in_data <= 8'hb5;
      11'd997  : in_data <= 8'h4e;
      11'd998  : in_data <= 8'h73;
      11'd999  : in_data <= 8'h6e;
      11'd1000 : in_data <= 8'hb5;
      11'd1001 : in_data <= 8'h61;
      11'd1002 : in_data <= 8'h3d;
      11'd1003 : in_data <= 8'h31;
      11'd1004 : in_data <= 8'h61;
      11'd1005 : in_data <= 8'h48;
      11'd1006 : in_data <= 8'h13;
      11'd1007 : in_data <= 8'hb2;
      11'd1008 : in_data <= 8'hed;
      11'd1009 : in_data <= 8'h93;
      11'd1010 : in_data <= 8'h53;
      11'd1011 : in_data <= 8'h42;
      11'd1012 : in_data <= 8'h8a;
      11'd1013 : in_data <= 8'hf0;
      11'd1014 : in_data <= 8'hf4;
      11'd1015 : in_data <= 8'hab;
      11'd1016 : in_data <= 8'hce;
      11'd1017 : in_data <= 8'h28;
      11'd1018 : in_data <= 8'h2c;
      11'd1019 : in_data <= 8'ha9;
      11'd1020 : in_data <= 8'hc2;
      11'd1021 : in_data <= 8'h34;
      11'd1022 : in_data <= 8'h30;
      11'd1023 : in_data <= 8'h03;
      11'd1024 : in_data <= 8'h7d;
      11'd1025 : in_data <= 8'h6b;
      11'd1026 : in_data <= 8'h33;
      11'd1027 : in_data <= 8'h6e;
      11'd1028 : in_data <= 8'h01;
      11'd1029 : in_data <= 8'h4b;
      11'd1030 : in_data <= 8'he6;
      11'd1031 : in_data <= 8'hab;
      11'd1032 : in_data <= 8'h6c;
      11'd1033 : in_data <= 8'h6a;
      11'd1034 : in_data <= 8'hca;
      11'd1035 : in_data <= 8'h57;
      11'd1036 : in_data <= 8'h5b;
      11'd1037 : in_data <= 8'h5f;
      11'd1038 : in_data <= 8'h0e;
      11'd1039 : in_data <= 8'hdf;
      11'd1040 : in_data <= 8'h35;
      11'd1041 : in_data <= 8'h9e;
      11'd1042 : in_data <= 8'h65;
      11'd1043 : in_data <= 8'h50;
      11'd1044 : in_data <= 8'hb6;
      11'd1045 : in_data <= 8'h4a;
      11'd1046 : in_data <= 8'he8;
      11'd1047 : in_data <= 8'hab;
      11'd1048 : in_data <= 8'h9d;
      11'd1049 : in_data <= 8'hbc;
      11'd1050 : in_data <= 8'h23;
      11'd1051 : in_data <= 8'h01;
      11'd1052 : in_data <= 8'h7d;
      11'd1053 : in_data <= 8'h71;
      11'd1054 : in_data <= 8'ha8;
      11'd1055 : in_data <= 8'h58;
      11'd1056 : in_data <= 8'hcc;
      11'd1057 : in_data <= 8'h6b;
      11'd1058 : in_data <= 8'ha4;
      11'd1059 : in_data <= 8'hf6;
      11'd1060 : in_data <= 8'h01;
      11'd1061 : in_data <= 8'h74;
      11'd1062 : in_data <= 8'h57;
      11'd1063 : in_data <= 8'heb;
      11'd1064 : in_data <= 8'hc3;
      11'd1065 : in_data <= 8'h7b;
      11'd1066 : in_data <= 8'hf8;
      11'd1067 : in_data <= 8'h4e;
      11'd1068 : in_data <= 8'h80;
      11'd1069 : in_data <= 8'h4d;
      11'd1070 : in_data <= 8'h1f;
      11'd1071 : in_data <= 8'h68;
      11'd1072 : in_data <= 8'hb6;
      11'd1073 : in_data <= 8'h71;
      11'd1074 : in_data <= 8'h5f;
      11'd1075 : in_data <= 8'h1d;
      11'd1076 : in_data <= 8'h22;
      11'd1077 : in_data <= 8'h33;
      11'd1078 : in_data <= 8'hcd;
      11'd1079 : in_data <= 8'hb4;
      11'd1080 : in_data <= 8'hc0;
      11'd1081 : in_data <= 8'hcf;
      11'd1082 : in_data <= 8'h0f;
      11'd1083 : in_data <= 8'hff;
      11'd1084 : in_data <= 8'ha5;
      11'd1085 : in_data <= 8'h82;
      11'd1086 : in_data <= 8'h78;
      11'd1087 : in_data <= 8'hcd;
      11'd1088 : in_data <= 8'ha7;
      11'd1089 : in_data <= 8'h9b;
      11'd1090 : in_data <= 8'h96;
      11'd1091 : in_data <= 8'h7c;
      11'd1092 : in_data <= 8'h7c;
      11'd1093 : in_data <= 8'h3d;
      11'd1094 : in_data <= 8'hd0;
      11'd1095 : in_data <= 8'h4d;
      11'd1096 : in_data <= 8'h20;
      11'd1097 : in_data <= 8'he0;
      11'd1098 : in_data <= 8'hc4;
      11'd1099 : in_data <= 8'h5c;
      11'd1100 : in_data <= 8'hf7;
      11'd1101 : in_data <= 8'h96;
      11'd1102 : in_data <= 8'h35;
      11'd1103 : in_data <= 8'hc7;
      11'd1104 : in_data <= 8'h58;
      11'd1105 : in_data <= 8'h6a;
      11'd1106 : in_data <= 8'ha0;
      11'd1107 : in_data <= 8'h3b;
      11'd1108 : in_data <= 8'ha0;
      11'd1109 : in_data <= 8'h03;
      11'd1110 : in_data <= 8'h70;
      11'd1111 : in_data <= 8'h80;
      11'd1112 : in_data <= 8'h3f;
      11'd1113 : in_data <= 8'h38;
      11'd1114 : in_data <= 8'h65;
      11'd1115 : in_data <= 8'h3b;
      11'd1116 : in_data <= 8'h39;
      11'd1117 : in_data <= 8'hbb;
      11'd1118 : in_data <= 8'hdd;
      11'd1119 : in_data <= 8'h40;
      11'd1120 : in_data <= 8'h43;
      11'd1121 : in_data <= 8'h9c;
      11'd1122 : in_data <= 8'h76;
      11'd1123 : in_data <= 8'h02;
      11'd1124 : in_data <= 8'h4d;
      11'd1125 : in_data <= 8'h18;
      11'd1126 : in_data <= 8'h16;
      11'd1127 : in_data <= 8'h75;
      11'd1128 : in_data <= 8'h78;
      11'd1129 : in_data <= 8'ha5;
      11'd1130 : in_data <= 8'hd4;
      11'd1131 : in_data <= 8'h27;
      11'd1132 : in_data <= 8'h3c;
      11'd1133 : in_data <= 8'hde;
      11'd1134 : in_data <= 8'hf9;
      11'd1135 : in_data <= 8'h7d;
      11'd1136 : in_data <= 8'he1;
      11'd1137 : in_data <= 8'hc9;
      11'd1138 : in_data <= 8'hb0;
      11'd1139 : in_data <= 8'h6e;
      11'd1140 : in_data <= 8'ha3;
      11'd1141 : in_data <= 8'h17;
      11'd1142 : in_data <= 8'h24;
      11'd1143 : in_data <= 8'hda;
      11'd1144 : in_data <= 8'h6f;
      11'd1145 : in_data <= 8'hbb;
      11'd1146 : in_data <= 8'hd8;
      11'd1147 : in_data <= 8'h2a;
      11'd1148 : in_data <= 8'had;
      11'd1149 : in_data <= 8'h0d;
      11'd1150 : in_data <= 8'h05;
      11'd1151 : in_data <= 8'h0d;
      11'd1152 : in_data <= 8'h91;
      11'd1153 : in_data <= 8'h65;
      11'd1154 : in_data <= 8'h75;
      11'd1155 : in_data <= 8'h1e;
      11'd1156 : in_data <= 8'h81;
      11'd1157 : in_data <= 8'h29;
      11'd1158 : in_data <= 8'h47;
      11'd1159 : in_data <= 8'h92;
      11'd1160 : in_data <= 8'h8c;
      11'd1161 : in_data <= 8'h94;
      11'd1162 : in_data <= 8'hc8;
      11'd1163 : in_data <= 8'h10;
      11'd1164 : in_data <= 8'h92;
      11'd1165 : in_data <= 8'hcf;
      11'd1166 : in_data <= 8'h5b;
      11'd1167 : in_data <= 8'hbf;
      11'd1168 : in_data <= 8'h81;
      11'd1169 : in_data <= 8'had;
      11'd1170 : in_data <= 8'hc6;
      11'd1171 : in_data <= 8'h87;
      11'd1172 : in_data <= 8'h74;
      11'd1173 : in_data <= 8'hfb;
      11'd1174 : in_data <= 8'h69;
      11'd1175 : in_data <= 8'h76;
      11'd1176 : in_data <= 8'h02;
      11'd1177 : in_data <= 8'hcc;
      11'd1178 : in_data <= 8'h52;
      11'd1179 : in_data <= 8'hbc;
      11'd1180 : in_data <= 8'h9e;
      11'd1181 : in_data <= 8'h1a;
      11'd1182 : in_data <= 8'hc7;
      11'd1183 : in_data <= 8'hfa;
      11'd1184 : in_data <= 8'h30;
      11'd1185 : in_data <= 8'h9e;
      11'd1186 : in_data <= 8'hb5;
      11'd1187 : in_data <= 8'hd2;
      11'd1188 : in_data <= 8'hb9;
      11'd1189 : in_data <= 8'h75;
      11'd1190 : in_data <= 8'he0;
      11'd1191 : in_data <= 8'hcb;
      11'd1192 : in_data <= 8'h0c;
      11'd1193 : in_data <= 8'ha7;
      11'd1194 : in_data <= 8'h93;
      11'd1195 : in_data <= 8'h20;
      11'd1196 : in_data <= 8'h06;
      11'd1197 : in_data <= 8'h1b;
      11'd1198 : in_data <= 8'h88;
      11'd1199 : in_data <= 8'h37;
      11'd1200 : in_data <= 8'h7a;
      11'd1201 : in_data <= 8'h47;
      11'd1202 : in_data <= 8'h57;
      11'd1203 : in_data <= 8'hcf;
      11'd1204 : in_data <= 8'h3a;
      11'd1205 : in_data <= 8'h26;
      11'd1206 : in_data <= 8'h2e;
      11'd1207 : in_data <= 8'h74;
      11'd1208 : in_data <= 8'h3d;
      11'd1209 : in_data <= 8'h6a;
      11'd1210 : in_data <= 8'h7b;
      11'd1211 : in_data <= 8'h10;
      11'd1212 : in_data <= 8'h3e;
      11'd1213 : in_data <= 8'h68;
      11'd1214 : in_data <= 8'h56;
      11'd1215 : in_data <= 8'h18;
      11'd1216 : in_data <= 8'h55;
      11'd1217 : in_data <= 8'h70;
      11'd1218 : in_data <= 8'h73;
      11'd1219 : in_data <= 8'hcb;
      11'd1220 : in_data <= 8'hc3;
      11'd1221 : in_data <= 8'h27;
      11'd1222 : in_data <= 8'h1e;
      11'd1223 : in_data <= 8'h48;
      11'd1224 : in_data <= 8'h68;
      11'd1225 : in_data <= 8'hc5;
      11'd1226 : in_data <= 8'h59;
      11'd1227 : in_data <= 8'h28;
      11'd1228 : in_data <= 8'hbb;
      11'd1229 : in_data <= 8'hcc;
      11'd1230 : in_data <= 8'h0b;
      11'd1231 : in_data <= 8'h5b;
      11'd1232 : in_data <= 8'h24;
      11'd1233 : in_data <= 8'hc1;
      11'd1234 : in_data <= 8'h2d;
      11'd1235 : in_data <= 8'h87;
      11'd1236 : in_data <= 8'h79;
      11'd1237 : in_data <= 8'h19;
      11'd1238 : in_data <= 8'h50;
      11'd1239 : in_data <= 8'hdf;
      11'd1240 : in_data <= 8'h94;
      11'd1241 : in_data <= 8'hbd;
      11'd1242 : in_data <= 8'h12;
      11'd1243 : in_data <= 8'h22;
      11'd1244 : in_data <= 8'hdb;
      11'd1245 : in_data <= 8'h5f;
      11'd1246 : in_data <= 8'he1;
      11'd1247 : in_data <= 8'h1f;
      11'd1248 : in_data <= 8'hce;
      11'd1249 : in_data <= 8'h72;
      11'd1250 : in_data <= 8'h98;
      11'd1251 : in_data <= 8'hc0;
      11'd1252 : in_data <= 8'h08;
      11'd1253 : in_data <= 8'h25;
      11'd1254 : in_data <= 8'h34;
      11'd1255 : in_data <= 8'h86;
      11'd1256 : in_data <= 8'h91;
      11'd1257 : in_data <= 8'hdb;
      11'd1258 : in_data <= 8'hb4;
      11'd1259 : in_data <= 8'h46;
      11'd1260 : in_data <= 8'ha6;
      11'd1261 : in_data <= 8'h98;
      11'd1262 : in_data <= 8'h33;
      11'd1263 : in_data <= 8'h9d;
      11'd1264 : in_data <= 8'hde;
      11'd1265 : in_data <= 8'h79;
      11'd1266 : in_data <= 8'h63;
      11'd1267 : in_data <= 8'hef;
      11'd1268 : in_data <= 8'h3e;
      11'd1269 : in_data <= 8'h9f;
      11'd1270 : in_data <= 8'hb4;
      11'd1271 : in_data <= 8'h8d;
      11'd1272 : in_data <= 8'hbe;
      11'd1273 : in_data <= 8'h4b;
      11'd1274 : in_data <= 8'hcc;
      11'd1275 : in_data <= 8'h93;
      11'd1276 : in_data <= 8'hb6;
      11'd1277 : in_data <= 8'h51;
      11'd1278 : in_data <= 8'h28;
      11'd1279 : in_data <= 8'h43;
      11'd1280 : in_data <= 8'h57;
      11'd1281 : in_data <= 8'hb2;
      11'd1282 : in_data <= 8'h72;
      11'd1283 : in_data <= 8'ha5;
      11'd1284 : in_data <= 8'h1b;
      11'd1285 : in_data <= 8'hd7;
      11'd1286 : in_data <= 8'h98;
      11'd1287 : in_data <= 8'h97;
      11'd1288 : in_data <= 8'h0d;
      11'd1289 : in_data <= 8'hba;
      11'd1290 : in_data <= 8'h15;
      11'd1291 : in_data <= 8'h6f;
      11'd1292 : in_data <= 8'h7b;
      11'd1293 : in_data <= 8'had;
      11'd1294 : in_data <= 8'h6c;
      11'd1295 : in_data <= 8'hfc;
      11'd1296 : in_data <= 8'h5e;
      11'd1297 : in_data <= 8'h9f;
      11'd1298 : in_data <= 8'hd1;
      11'd1299 : in_data <= 8'h1f;
      11'd1300 : in_data <= 8'h8e;
      11'd1301 : in_data <= 8'h94;
      11'd1302 : in_data <= 8'ha4;
      11'd1303 : in_data <= 8'h45;
      11'd1304 : in_data <= 8'h10;
      11'd1305 : in_data <= 8'h75;
      11'd1306 : in_data <= 8'h0d;
      11'd1307 : in_data <= 8'hb4;
      11'd1308 : in_data <= 8'h63;
      11'd1309 : in_data <= 8'hde;
      11'd1310 : in_data <= 8'hc6;
      11'd1311 : in_data <= 8'h25;
      11'd1312 : in_data <= 8'h94;
      11'd1313 : in_data <= 8'h07;
      11'd1314 : in_data <= 8'h59;
      11'd1315 : in_data <= 8'h59;
      11'd1316 : in_data <= 8'h7c;
      11'd1317 : in_data <= 8'hee;
      11'd1318 : in_data <= 8'h24;
      11'd1319 : in_data <= 8'h53;
      11'd1320 : in_data <= 8'h83;
      11'd1321 : in_data <= 8'hda;
      11'd1322 : in_data <= 8'ha8;
      11'd1323 : in_data <= 8'hc1;
      11'd1324 : in_data <= 8'h06;
      11'd1325 : in_data <= 8'h9e;
      11'd1326 : in_data <= 8'ha1;
      11'd1327 : in_data <= 8'hb4;
      11'd1328 : in_data <= 8'h38;
      11'd1329 : in_data <= 8'h1d;
      11'd1330 : in_data <= 8'he6;
      11'd1331 : in_data <= 8'hd5;
      11'd1332 : in_data <= 8'h74;
      11'd1333 : in_data <= 8'h52;
      11'd1334 : in_data <= 8'hf9;
      11'd1335 : in_data <= 8'h25;
      11'd1336 : in_data <= 8'h69;
      11'd1337 : in_data <= 8'h44;
      11'd1338 : in_data <= 8'h53;
      11'd1339 : in_data <= 8'he2;
      11'd1340 : in_data <= 8'h35;
      11'd1341 : in_data <= 8'h6d;
      11'd1342 : in_data <= 8'h09;
      11'd1343 : in_data <= 8'h62;
      11'd1344 : in_data <= 8'h15;
      11'd1345 : in_data <= 8'h64;
      11'd1346 : in_data <= 8'h38;
      11'd1347 : in_data <= 8'h8b;
      11'd1348 : in_data <= 8'h3f;
      11'd1349 : in_data <= 8'h17;
      11'd1350 : in_data <= 8'hd1;
      11'd1351 : in_data <= 8'hcc;
      11'd1352 : in_data <= 8'hb8;
      11'd1353 : in_data <= 8'h77;
      11'd1354 : in_data <= 8'h4a;
      11'd1355 : in_data <= 8'h22;
      11'd1356 : in_data <= 8'h51;
      11'd1357 : in_data <= 8'hf5;
      11'd1358 : in_data <= 8'hba;
      11'd1359 : in_data <= 8'h57;
      11'd1360 : in_data <= 8'hc4;
      11'd1361 : in_data <= 8'hce;
      11'd1362 : in_data <= 8'h20;
      11'd1363 : in_data <= 8'hcf;
      11'd1364 : in_data <= 8'h98;
      11'd1365 : in_data <= 8'h32;
      11'd1366 : in_data <= 8'h97;
      11'd1367 : in_data <= 8'h0a;
      11'd1368 : in_data <= 8'hbe;
      11'd1369 : in_data <= 8'h30;
      11'd1370 : in_data <= 8'hf3;
      11'd1371 : in_data <= 8'h1f;
      11'd1372 : in_data <= 8'he6;
      11'd1373 : in_data <= 8'h55;
      11'd1374 : in_data <= 8'h1e;
      11'd1375 : in_data <= 8'ha8;
      11'd1376 : in_data <= 8'h42;
      11'd1377 : in_data <= 8'hd8;
      11'd1378 : in_data <= 8'h3d;
      11'd1379 : in_data <= 8'hc2;
      11'd1380 : in_data <= 8'hb3;
      11'd1381 : in_data <= 8'hf5;
      11'd1382 : in_data <= 8'heb;
      11'd1383 : in_data <= 8'hb5;
      11'd1384 : in_data <= 8'hdb;
      11'd1385 : in_data <= 8'hea;
      11'd1386 : in_data <= 8'h6f;
      11'd1387 : in_data <= 8'h7a;
      11'd1388 : in_data <= 8'hb9;
      11'd1389 : in_data <= 8'h85;
      11'd1390 : in_data <= 8'h40;
      11'd1391 : in_data <= 8'h2b;
      11'd1392 : in_data <= 8'h05;
      11'd1393 : in_data <= 8'ha5;
      11'd1394 : in_data <= 8'h28;
      11'd1395 : in_data <= 8'h90;
      11'd1396 : in_data <= 8'he6;
      11'd1397 : in_data <= 8'h26;
      11'd1398 : in_data <= 8'h83;
      11'd1399 : in_data <= 8'h14;
      11'd1400 : in_data <= 8'h30;
      11'd1401 : in_data <= 8'hac;
      11'd1402 : in_data <= 8'hd5;
      11'd1403 : in_data <= 8'hae;
      11'd1404 : in_data <= 8'h68;
      11'd1405 : in_data <= 8'hb6;
      11'd1406 : in_data <= 8'h67;
      11'd1407 : in_data <= 8'h2e;
      11'd1408 : in_data <= 8'h09;
      11'd1409 : in_data <= 8'hed;
      11'd1410 : in_data <= 8'h35;
      11'd1411 : in_data <= 8'h4a;
      11'd1412 : in_data <= 8'hef;
      11'd1413 : in_data <= 8'h48;
      11'd1414 : in_data <= 8'h90;
      11'd1415 : in_data <= 8'h57;
      11'd1416 : in_data <= 8'h9f;
      11'd1417 : in_data <= 8'h41;
      11'd1418 : in_data <= 8'h7e;
      11'd1419 : in_data <= 8'h80;
      11'd1420 : in_data <= 8'h43;
      11'd1421 : in_data <= 8'h6f;
      11'd1422 : in_data <= 8'hf5;
      11'd1423 : in_data <= 8'hf7;
      11'd1424 : in_data <= 8'h88;
      11'd1425 : in_data <= 8'hb1;
      11'd1426 : in_data <= 8'ha9;
      11'd1427 : in_data <= 8'h16;
      11'd1428 : in_data <= 8'h0a;
      11'd1429 : in_data <= 8'h50;
      11'd1430 : in_data <= 8'h24;
      11'd1431 : in_data <= 8'hf3;
      11'd1432 : in_data <= 8'h55;
      11'd1433 : in_data <= 8'hfc;
      11'd1434 : in_data <= 8'hb6;
      11'd1435 : in_data <= 8'hf5;
      11'd1436 : in_data <= 8'hc8;
      11'd1437 : in_data <= 8'h7b;
      11'd1438 : in_data <= 8'hea;
      11'd1439 : in_data <= 8'hef;
      11'd1440 : in_data <= 8'h23;
      11'd1441 : in_data <= 8'h87;
      11'd1442 : in_data <= 8'h25;
      11'd1443 : in_data <= 8'h08;
      11'd1444 : in_data <= 8'h11;
      11'd1445 : in_data <= 8'had;
      11'd1446 : in_data <= 8'h1c;
      11'd1447 : in_data <= 8'ha6;
      11'd1448 : in_data <= 8'he8;
      11'd1449 : in_data <= 8'h1a;
      11'd1450 : in_data <= 8'h29;
      11'd1451 : in_data <= 8'hc0;
      11'd1452 : in_data <= 8'hae;
      11'd1453 : in_data <= 8'heb;
      11'd1454 : in_data <= 8'h13;
      11'd1455 : in_data <= 8'h09;
      11'd1456 : in_data <= 8'h45;
      11'd1457 : in_data <= 8'h63;
      11'd1458 : in_data <= 8'h3a;
      11'd1459 : in_data <= 8'h3c;
      11'd1460 : in_data <= 8'hef;
      11'd1461 : in_data <= 8'hd7;
      11'd1462 : in_data <= 8'h8b;
      11'd1463 : in_data <= 8'hf6;
      11'd1464 : in_data <= 8'ha4;
      11'd1465 : in_data <= 8'h03;
      11'd1466 : in_data <= 8'h77;
      11'd1467 : in_data <= 8'hb4;
      11'd1468 : in_data <= 8'h33;
      11'd1469 : in_data <= 8'hbc;
      11'd1470 : in_data <= 8'h59;
      11'd1471 : in_data <= 8'hff;
      11'd1472 : in_data <= 8'h4f;
      11'd1473 : in_data <= 8'hac;
      11'd1474 : in_data <= 8'h60;
      11'd1475 : in_data <= 8'h33;
      11'd1476 : in_data <= 8'h42;
      11'd1477 : in_data <= 8'h78;
      11'd1478 : in_data <= 8'h35;
      11'd1479 : in_data <= 8'hfe;
      11'd1480 : in_data <= 8'h62;
      11'd1481 : in_data <= 8'hd3;
      11'd1482 : in_data <= 8'hb0;
      11'd1483 : in_data <= 8'h5f;
      11'd1484 : in_data <= 8'hcb;
      11'd1485 : in_data <= 8'h22;
      11'd1486 : in_data <= 8'h3d;
      11'd1487 : in_data <= 8'h40;
      11'd1488 : in_data <= 8'hfe;
      11'd1489 : in_data <= 8'h09;
      11'd1490 : in_data <= 8'h49;
      11'd1491 : in_data <= 8'h5d;
      11'd1492 : in_data <= 8'he3;
      11'd1493 : in_data <= 8'h1b;
      11'd1494 : in_data <= 8'hbc;
      11'd1495 : in_data <= 8'h0c;
      11'd1496 : in_data <= 8'hb3;
      11'd1497 : in_data <= 8'h0a;
      11'd1498 : in_data <= 8'h97;
      11'd1499 : in_data <= 8'hb2;
      11'd1500 : in_data <= 8'h34;
      11'd1501 : in_data <= 8'hee;
      11'd1502 : in_data <= 8'h43;
      11'd1503 : in_data <= 8'h6c;
      11'd1504 : in_data <= 8'h87;
      11'd1505 : in_data <= 8'h3f;
      11'd1506 : in_data <= 8'he3;
      11'd1507 : in_data <= 8'h2e;
      11'd1508 : in_data <= 8'hcb;
      11'd1509 : in_data <= 8'he4;
      11'd1510 : in_data <= 8'h59;
      11'd1511 : in_data <= 8'h2b;
      11'd1512 : in_data <= 8'hd7;
      11'd1513 : in_data <= 8'hb8;
      11'd1514 : in_data <= 8'h36;
      11'd1515 : in_data <= 8'hb3;
      11'd1516 : in_data <= 8'h8d;
      11'd1517 : in_data <= 8'hc3;
      11'd1518 : in_data <= 8'hbe;
      11'd1519 : in_data <= 8'h8c;
      11'd1520 : in_data <= 8'hc7;
      11'd1521 : in_data <= 8'h98;
      11'd1522 : in_data <= 8'h96;
      11'd1523 : in_data <= 8'h88;
      11'd1524 : in_data <= 8'h5f;
      11'd1525 : in_data <= 8'hbc;
      11'd1526 : in_data <= 8'h16;
      11'd1527 : in_data <= 8'hcb;
      11'd1528 : in_data <= 8'he7;
      11'd1529 : in_data <= 8'he7;
      11'd1530 : in_data <= 8'h58;
      11'd1531 : in_data <= 8'h45;
      11'd1532 : in_data <= 8'hfc;
      11'd1533 : in_data <= 8'h7a;
      11'd1534 : in_data <= 8'h12;
      11'd1535 : in_data <= 8'h9b;
      11'd1536 : in_data <= 8'h21;
      11'd1537 : in_data <= 8'h2b;
      11'd1538 : in_data <= 8'had;
      11'd1539 : in_data <= 8'hc5;
      11'd1540 : in_data <= 8'h22;
      11'd1541 : in_data <= 8'hf6;
      11'd1542 : in_data <= 8'h47;
      11'd1543 : in_data <= 8'hb5;
      11'd1544 : in_data <= 8'h37;
      11'd1545 : in_data <= 8'hdc;
      11'd1546 : in_data <= 8'h75;
      11'd1547 : in_data <= 8'he7;
      11'd1548 : in_data <= 8'h51;
      11'd1549 : in_data <= 8'hef;
      11'd1550 : in_data <= 8'h1f;
      11'd1551 : in_data <= 8'h14;
      11'd1552 : in_data <= 8'h41;
      11'd1553 : in_data <= 8'hca;
      11'd1554 : in_data <= 8'hab;
      11'd1555 : in_data <= 8'h23;
      11'd1556 : in_data <= 8'hc4;
      11'd1557 : in_data <= 8'h23;
      11'd1558 : in_data <= 8'h33;
      11'd1559 : in_data <= 8'h29;
      11'd1560 : in_data <= 8'h12;
      11'd1561 : in_data <= 8'h75;
      11'd1562 : in_data <= 8'hfd;
      11'd1563 : in_data <= 8'h03;
      11'd1564 : in_data <= 8'hb7;
      11'd1565 : in_data <= 8'ha4;
      11'd1566 : in_data <= 8'hb4;
      11'd1567 : in_data <= 8'hb4;
      11'd1568 : in_data <= 8'h96;
      11'd1569 : in_data <= 8'h45;
      11'd1570 : in_data <= 8'he1;
      11'd1571 : in_data <= 8'hac;
      11'd1572 : in_data <= 8'h0f;
      11'd1573 : in_data <= 8'he5;
      11'd1574 : in_data <= 8'h84;
      11'd1575 : in_data <= 8'h28;
      11'd1576 : in_data <= 8'h11;
      11'd1577 : in_data <= 8'h61;
      11'd1578 : in_data <= 8'hae;
      11'd1579 : in_data <= 8'h92;
      11'd1580 : in_data <= 8'h4a;
      11'd1581 : in_data <= 8'ha6;
      11'd1582 : in_data <= 8'h37;
      11'd1583 : in_data <= 8'h67;
      11'd1584 : in_data <= 8'h74;
      11'd1585 : in_data <= 8'h1c;
      11'd1586 : in_data <= 8'h32;
      11'd1587 : in_data <= 8'h33;
      11'd1588 : in_data <= 8'h51;
      11'd1589 : in_data <= 8'hde;
      11'd1590 : in_data <= 8'he4;
      11'd1591 : in_data <= 8'h7f;
      11'd1592 : in_data <= 8'hbe;
      11'd1593 : in_data <= 8'h14;
      11'd1594 : in_data <= 8'h2a;
      11'd1595 : in_data <= 8'ha2;
      11'd1596 : in_data <= 8'h66;
      11'd1597 : in_data <= 8'h4a;
      11'd1598 : in_data <= 8'h27;
      11'd1599 : in_data <= 8'hcd;
      11'd1600 : in_data <= 8'hda;
      11'd1601 : in_data <= 8'ha2;
      11'd1602 : in_data <= 8'hd6;
      11'd1603 : in_data <= 8'h0d;
      11'd1604 : in_data <= 8'hb8;
      11'd1605 : in_data <= 8'h35;
      11'd1606 : in_data <= 8'h74;
      11'd1607 : in_data <= 8'h47;
      11'd1608 : in_data <= 8'hc5;
      11'd1609 : in_data <= 8'h04;
      11'd1610 : in_data <= 8'h64;
      11'd1611 : in_data <= 8'hbf;
      11'd1612 : in_data <= 8'hfd;
      11'd1613 : in_data <= 8'h6e;
      11'd1614 : in_data <= 8'h11;
      11'd1615 : in_data <= 8'h1e;
      11'd1616 : in_data <= 8'h8d;
      11'd1617 : in_data <= 8'h38;
      11'd1618 : in_data <= 8'h25;
      11'd1619 : in_data <= 8'h7f;
      11'd1620 : in_data <= 8'h21;
      11'd1621 : in_data <= 8'h89;
      11'd1622 : in_data <= 8'had;
      11'd1623 : in_data <= 8'h64;
      11'd1624 : in_data <= 8'h1b;
      11'd1625 : in_data <= 8'hf8;
      11'd1626 : in_data <= 8'h1b;
      11'd1627 : in_data <= 8'hda;
      11'd1628 : in_data <= 8'h94;
      11'd1629 : in_data <= 8'h09;
      11'd1630 : in_data <= 8'h1d;
      11'd1631 : in_data <= 8'h49;
      11'd1632 : in_data <= 8'ha6;
      11'd1633 : in_data <= 8'h19;
      11'd1634 : in_data <= 8'h6e;
      11'd1635 : in_data <= 8'he3;
      11'd1636 : in_data <= 8'hda;
      11'd1637 : in_data <= 8'had;
      11'd1638 : in_data <= 8'hbc;
      11'd1639 : in_data <= 8'h5d;
      11'd1640 : in_data <= 8'h80;
      11'd1641 : in_data <= 8'h06;
      11'd1642 : in_data <= 8'h5c;
      11'd1643 : in_data <= 8'hcd;
      11'd1644 : in_data <= 8'h85;
      11'd1645 : in_data <= 8'h46;
      11'd1646 : in_data <= 8'h7e;
      11'd1647 : in_data <= 8'h82;
      11'd1648 : in_data <= 8'h4f;
      11'd1649 : in_data <= 8'ha8;
      11'd1650 : in_data <= 8'hac;
      11'd1651 : in_data <= 8'h89;
      11'd1652 : in_data <= 8'hbb;
      11'd1653 : in_data <= 8'h86;
      11'd1654 : in_data <= 8'h26;
      11'd1655 : in_data <= 8'ha1;
      11'd1656 : in_data <= 8'hdf;
      11'd1657 : in_data <= 8'hf0;
      11'd1658 : in_data <= 8'h89;
      11'd1659 : in_data <= 8'hc3;
      11'd1660 : in_data <= 8'hf9;
      11'd1661 : in_data <= 8'hbf;
      11'd1662 : in_data <= 8'h60;
      11'd1663 : in_data <= 8'h22;
      11'd1664 : in_data <= 8'h12;
      11'd1665 : in_data <= 8'hae;
      11'd1666 : in_data <= 8'h61;
      11'd1667 : in_data <= 8'h18;
      11'd1668 : in_data <= 8'h72;
      11'd1669 : in_data <= 8'h71;
      11'd1670 : in_data <= 8'h9e;
      11'd1671 : in_data <= 8'h95;
      11'd1672 : in_data <= 8'hcc;
      11'd1673 : in_data <= 8'hbd;
      11'd1674 : in_data <= 8'h01;
      11'd1675 : in_data <= 8'h6f;
      11'd1676 : in_data <= 8'h56;
      11'd1677 : in_data <= 8'h8c;
      11'd1678 : in_data <= 8'h95;
      11'd1679 : in_data <= 8'h11;
      11'd1680 : in_data <= 8'h77;
      11'd1681 : in_data <= 8'hf7;
      11'd1682 : in_data <= 8'hce;
      11'd1683 : in_data <= 8'h33;
      11'd1684 : in_data <= 8'h4e;
      11'd1685 : in_data <= 8'hde;
      11'd1686 : in_data <= 8'hd3;
      11'd1687 : in_data <= 8'hcc;
      11'd1688 : in_data <= 8'hab;
      11'd1689 : in_data <= 8'h2e;
      11'd1690 : in_data <= 8'hed;
      11'd1691 : in_data <= 8'h16;
      11'd1692 : in_data <= 8'hbc;
      11'd1693 : in_data <= 8'hc6;
      11'd1694 : in_data <= 8'hba;
      11'd1695 : in_data <= 8'h0a;
      11'd1696 : in_data <= 8'h49;
      11'd1697 : in_data <= 8'h08;
      11'd1698 : in_data <= 8'ha3;
      11'd1699 : in_data <= 8'h1d;
      11'd1700 : in_data <= 8'hfa;
      11'd1701 : in_data <= 8'ha2;
      11'd1702 : in_data <= 8'hcb;
      11'd1703 : in_data <= 8'hf2;
      11'd1704 : in_data <= 8'h96;
      11'd1705 : in_data <= 8'h1b;
      11'd1706 : in_data <= 8'hfc;
      11'd1707 : in_data <= 8'h65;
      11'd1708 : in_data <= 8'h09;
      11'd1709 : in_data <= 8'h6f;
      11'd1710 : in_data <= 8'ha4;
      11'd1711 : in_data <= 8'h33;
      11'd1712 : in_data <= 8'h0c;
      11'd1713 : in_data <= 8'h2d;
      11'd1714 : in_data <= 8'h01;
      11'd1715 : in_data <= 8'hd5;
      11'd1716 : in_data <= 8'h13;
      11'd1717 : in_data <= 8'h70;
      11'd1718 : in_data <= 8'h32;
      11'd1719 : in_data <= 8'he3;
      11'd1720 : in_data <= 8'h33;
      11'd1721 : in_data <= 8'h06;
      11'd1722 : in_data <= 8'he7;
      11'd1723 : in_data <= 8'h03;
      11'd1724 : in_data <= 8'hca;
      11'd1725 : in_data <= 8'h95;
      11'd1726 : in_data <= 8'h30;
      11'd1727 : in_data <= 8'h85;
      11'd1728 : in_data <= 8'ha0;
      11'd1729 : in_data <= 8'hb2;
      11'd1730 : in_data <= 8'h2c;
      11'd1731 : in_data <= 8'hbd;
      11'd1732 : in_data <= 8'ha7;
      11'd1733 : in_data <= 8'h25;
      11'd1734 : in_data <= 8'ha8;
      11'd1735 : in_data <= 8'h15;
      11'd1736 : in_data <= 8'h9b;
      11'd1737 : in_data <= 8'h62;
      11'd1738 : in_data <= 8'h8b;
      11'd1739 : in_data <= 8'h31;
      11'd1740 : in_data <= 8'ha6;
      11'd1741 : in_data <= 8'ha5;
      11'd1742 : in_data <= 8'h0e;
      11'd1743 : in_data <= 8'h4a;
      11'd1744 : in_data <= 8'h4a;
      11'd1745 : in_data <= 8'h56;
      11'd1746 : in_data <= 8'h20;
      11'd1747 : in_data <= 8'hf7;
      11'd1748 : in_data <= 8'h8f;
      11'd1749 : in_data <= 8'h19;
      11'd1750 : in_data <= 8'hd8;
      11'd1751 : in_data <= 8'h63;
      11'd1752 : in_data <= 8'h50;
      11'd1753 : in_data <= 8'hcd;
      11'd1754 : in_data <= 8'h38;
      11'd1755 : in_data <= 8'h73;
      11'd1756 : in_data <= 8'h1f;
      11'd1757 : in_data <= 8'hee;
      11'd1758 : in_data <= 8'ha5;
      11'd1759 : in_data <= 8'hb6;
      11'd1760 : in_data <= 8'h01;
      11'd1761 : in_data <= 8'hd6;
      11'd1762 : in_data <= 8'h44;
      11'd1763 : in_data <= 8'hd8;
      11'd1764 : in_data <= 8'h79;
      11'd1765 : in_data <= 8'hb2;
      11'd1766 : in_data <= 8'h3b;
      11'd1767 : in_data <= 8'hff;
      11'd1768 : in_data <= 8'h5a;
      11'd1769 : in_data <= 8'h2b;
      11'd1770 : in_data <= 8'hb6;
      11'd1771 : in_data <= 8'hcf;
      11'd1772 : in_data <= 8'h41;
      11'd1773 : in_data <= 8'h8d;
      11'd1774 : in_data <= 8'he2;
      11'd1775 : in_data <= 8'h4d;
      11'd1776 : in_data <= 8'h68;
      11'd1777 : in_data <= 8'h5c;
      11'd1778 : in_data <= 8'h3f;
      11'd1779 : in_data <= 8'hde;
      11'd1780 : in_data <= 8'h2a;
      11'd1781 : in_data <= 8'h67;
      11'd1782 : in_data <= 8'h7d;
      11'd1783 : in_data <= 8'h18;
      11'd1784 : in_data <= 8'h83;
      11'd1785 : in_data <= 8'h06;
      11'd1786 : in_data <= 8'h40;
      11'd1787 : in_data <= 8'h4d;
      11'd1788 : in_data <= 8'h57;
      11'd1789 : in_data <= 8'h3f;
      11'd1790 : in_data <= 8'hf9;
      11'd1791 : in_data <= 8'h28;
      11'd1792 : in_data <= 8'hda;
      11'd1793 : in_data <= 8'ha6;
      11'd1794 : in_data <= 8'ha6;
      11'd1795 : in_data <= 8'h75;
      11'd1796 : in_data <= 8'h57;
      11'd1797 : in_data <= 8'h0f;
      11'd1798 : in_data <= 8'h6c;
      11'd1799 : in_data <= 8'hc2;
      11'd1800 : in_data <= 8'hd0;
      11'd1801 : in_data <= 8'h59;
      11'd1802 : in_data <= 8'h8d;
      11'd1803 : in_data <= 8'hc2;
      11'd1804 : in_data <= 8'hf4;
      11'd1805 : in_data <= 8'hb5;
      11'd1806 : in_data <= 8'h9f;
      11'd1807 : in_data <= 8'h82;
      11'd1808 : in_data <= 8'hde;
      11'd1809 : in_data <= 8'h3d;
      11'd1810 : in_data <= 8'hac;
      11'd1811 : in_data <= 8'h31;
      11'd1812 : in_data <= 8'h4a;
      11'd1813 : in_data <= 8'h27;
      11'd1814 : in_data <= 8'h00;
      default: in_data <= 8'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      11'd0    : out_data_ref <= 14'h028c; // 'd652
      11'd1    : out_data_ref <= 14'h00d4; // 'd212
      11'd2    : out_data_ref <= 14'h047a; // 'd1146
      11'd3    : out_data_ref <= 14'h0826; // 'd2086
      11'd4    : out_data_ref <= 14'h015d; // 'd349
      11'd5    : out_data_ref <= 14'h09cc; // 'd2508
      11'd6    : out_data_ref <= 14'h0185; // 'd389
      11'd7    : out_data_ref <= 14'h0a33; // 'd2611
      11'd8    : out_data_ref <= 14'h0294; // 'd660
      11'd9    : out_data_ref <= 14'h01f7; // 'd503
      11'd10   : out_data_ref <= 14'h00f0; // 'd240
      11'd11   : out_data_ref <= 14'h06dd; // 'd1757
      11'd12   : out_data_ref <= 14'h0990; // 'd2448
      11'd13   : out_data_ref <= 14'h099b; // 'd2459
      11'd14   : out_data_ref <= 14'h0716; // 'd1814
      11'd15   : out_data_ref <= 14'h0038; // 'd56
      11'd16   : out_data_ref <= 14'h074b; // 'd1867
      11'd17   : out_data_ref <= 14'h053b; // 'd1339
      11'd18   : out_data_ref <= 14'h0770; // 'd1904
      11'd19   : out_data_ref <= 14'h0093; // 'd147
      11'd20   : out_data_ref <= 14'h06fd; // 'd1789
      11'd21   : out_data_ref <= 14'h03c4; // 'd964
      11'd22   : out_data_ref <= 14'h00b3; // 'd179
      11'd23   : out_data_ref <= 14'h09b1; // 'd2481
      11'd24   : out_data_ref <= 14'h05e1; // 'd1505
      11'd25   : out_data_ref <= 14'h09c7; // 'd2503
      11'd26   : out_data_ref <= 14'h03ac; // 'd940
      11'd27   : out_data_ref <= 14'h0603; // 'd1539
      11'd28   : out_data_ref <= 14'h00fe; // 'd254
      11'd29   : out_data_ref <= 14'h0730; // 'd1840
      11'd30   : out_data_ref <= 14'h05f3; // 'd1523
      11'd31   : out_data_ref <= 14'h02d5; // 'd725
      11'd32   : out_data_ref <= 14'h0295; // 'd661
      11'd33   : out_data_ref <= 14'h0370; // 'd880
      11'd34   : out_data_ref <= 14'h0839; // 'd2105
      11'd35   : out_data_ref <= 14'h09bf; // 'd2495
      11'd36   : out_data_ref <= 14'h07cc; // 'd1996
      11'd37   : out_data_ref <= 14'h04ad; // 'd1197
      11'd38   : out_data_ref <= 14'h0956; // 'd2390
      11'd39   : out_data_ref <= 14'h0676; // 'd1654
      11'd40   : out_data_ref <= 14'h0343; // 'd835
      11'd41   : out_data_ref <= 14'h00df; // 'd223
      11'd42   : out_data_ref <= 14'h07f4; // 'd2036
      11'd43   : out_data_ref <= 14'h0807; // 'd2055
      11'd44   : out_data_ref <= 14'h0055; // 'd85
      11'd45   : out_data_ref <= 14'h047b; // 'd1147
      11'd46   : out_data_ref <= 14'h05c9; // 'd1481
      11'd47   : out_data_ref <= 14'h085d; // 'd2141
      11'd48   : out_data_ref <= 14'h04a6; // 'd1190
      11'd49   : out_data_ref <= 14'h0155; // 'd341
      11'd50   : out_data_ref <= 14'h05f6; // 'd1526
      11'd51   : out_data_ref <= 14'h079b; // 'd1947
      11'd52   : out_data_ref <= 14'h02aa; // 'd682
      11'd53   : out_data_ref <= 14'h0219; // 'd537
      11'd54   : out_data_ref <= 14'h02fe; // 'd766
      11'd55   : out_data_ref <= 14'h0006; // 'd6
      11'd56   : out_data_ref <= 14'h095c; // 'd2396
      11'd57   : out_data_ref <= 14'h075c; // 'd1884
      11'd58   : out_data_ref <= 14'h03ed; // 'd1005
      11'd59   : out_data_ref <= 14'h014f; // 'd335
      11'd60   : out_data_ref <= 14'h09e2; // 'd2530
      11'd61   : out_data_ref <= 14'h0a26; // 'd2598
      11'd62   : out_data_ref <= 14'h053d; // 'd1341
      11'd63   : out_data_ref <= 14'h05fd; // 'd1533
      11'd64   : out_data_ref <= 14'h09c4; // 'd2500
      11'd65   : out_data_ref <= 14'h0784; // 'd1924
      11'd66   : out_data_ref <= 14'h06e3; // 'd1763
      11'd67   : out_data_ref <= 14'h0687; // 'd1671
      11'd68   : out_data_ref <= 14'h043b; // 'd1083
      11'd69   : out_data_ref <= 14'h071b; // 'd1819
      11'd70   : out_data_ref <= 14'h00e7; // 'd231
      11'd71   : out_data_ref <= 14'h080c; // 'd2060
      11'd72   : out_data_ref <= 14'h0873; // 'd2163
      11'd73   : out_data_ref <= 14'h07d1; // 'd2001
      11'd74   : out_data_ref <= 14'h0997; // 'd2455
      11'd75   : out_data_ref <= 14'h093b; // 'd2363
      11'd76   : out_data_ref <= 14'h083b; // 'd2107
      11'd77   : out_data_ref <= 14'h012e; // 'd302
      11'd78   : out_data_ref <= 14'h0522; // 'd1314
      11'd79   : out_data_ref <= 14'h01a2; // 'd418
      11'd80   : out_data_ref <= 14'h0681; // 'd1665
      11'd81   : out_data_ref <= 14'h0893; // 'd2195
      11'd82   : out_data_ref <= 14'h0692; // 'd1682
      11'd83   : out_data_ref <= 14'h0918; // 'd2328
      11'd84   : out_data_ref <= 14'h0a0f; // 'd2575
      11'd85   : out_data_ref <= 14'h085b; // 'd2139
      11'd86   : out_data_ref <= 14'h040a; // 'd1034
      11'd87   : out_data_ref <= 14'h0359; // 'd857
      11'd88   : out_data_ref <= 14'h0618; // 'd1560
      11'd89   : out_data_ref <= 14'h0090; // 'd144
      11'd90   : out_data_ref <= 14'h09ed; // 'd2541
      11'd91   : out_data_ref <= 14'h092c; // 'd2348
      11'd92   : out_data_ref <= 14'h0838; // 'd2104
      11'd93   : out_data_ref <= 14'h0453; // 'd1107
      11'd94   : out_data_ref <= 14'h0849; // 'd2121
      11'd95   : out_data_ref <= 14'h0166; // 'd358
      11'd96   : out_data_ref <= 14'h0824; // 'd2084
      11'd97   : out_data_ref <= 14'h07a7; // 'd1959
      11'd98   : out_data_ref <= 14'h06c3; // 'd1731
      11'd99   : out_data_ref <= 14'h06a6; // 'd1702
      11'd100  : out_data_ref <= 14'h020c; // 'd524
      11'd101  : out_data_ref <= 14'h0105; // 'd261
      11'd102  : out_data_ref <= 14'h0851; // 'd2129
      11'd103  : out_data_ref <= 14'h0622; // 'd1570
      11'd104  : out_data_ref <= 14'h010b; // 'd267
      11'd105  : out_data_ref <= 14'h00fb; // 'd251
      11'd106  : out_data_ref <= 14'h0503; // 'd1283
      11'd107  : out_data_ref <= 14'h0340; // 'd832
      11'd108  : out_data_ref <= 14'h027d; // 'd637
      11'd109  : out_data_ref <= 14'h03b5; // 'd949
      11'd110  : out_data_ref <= 14'h0573; // 'd1395
      11'd111  : out_data_ref <= 14'h07c0; // 'd1984
      11'd112  : out_data_ref <= 14'h08e8; // 'd2280
      11'd113  : out_data_ref <= 14'h0710; // 'd1808
      11'd114  : out_data_ref <= 14'h062d; // 'd1581
      11'd115  : out_data_ref <= 14'h0173; // 'd371
      11'd116  : out_data_ref <= 14'h0614; // 'd1556
      11'd117  : out_data_ref <= 14'h062b; // 'd1579
      11'd118  : out_data_ref <= 14'h093d; // 'd2365
      11'd119  : out_data_ref <= 14'h0460; // 'd1120
      11'd120  : out_data_ref <= 14'h0776; // 'd1910
      11'd121  : out_data_ref <= 14'h03d7; // 'd983
      11'd122  : out_data_ref <= 14'h0a2e; // 'd2606
      11'd123  : out_data_ref <= 14'h0857; // 'd2135
      11'd124  : out_data_ref <= 14'h09bd; // 'd2493
      11'd125  : out_data_ref <= 14'h0254; // 'd596
      11'd126  : out_data_ref <= 14'h0280; // 'd640
      11'd127  : out_data_ref <= 14'h069e; // 'd1694
      11'd128  : out_data_ref <= 14'h0601; // 'd1537
      11'd129  : out_data_ref <= 14'h0083; // 'd131
      11'd130  : out_data_ref <= 14'h06bc; // 'd1724
      11'd131  : out_data_ref <= 14'h09ae; // 'd2478
      11'd132  : out_data_ref <= 14'h02fa; // 'd762
      11'd133  : out_data_ref <= 14'h03b5; // 'd949
      11'd134  : out_data_ref <= 14'h00d1; // 'd209
      11'd135  : out_data_ref <= 14'h0541; // 'd1345
      11'd136  : out_data_ref <= 14'h00c2; // 'd194
      11'd137  : out_data_ref <= 14'h00fd; // 'd253
      11'd138  : out_data_ref <= 14'h0662; // 'd1634
      11'd139  : out_data_ref <= 14'h015d; // 'd349
      11'd140  : out_data_ref <= 14'h0097; // 'd151
      11'd141  : out_data_ref <= 14'h0548; // 'd1352
      11'd142  : out_data_ref <= 14'h0560; // 'd1376
      11'd143  : out_data_ref <= 14'h0a10; // 'd2576
      11'd144  : out_data_ref <= 14'h0677; // 'd1655
      11'd145  : out_data_ref <= 14'h0704; // 'd1796
      11'd146  : out_data_ref <= 14'h0751; // 'd1873
      11'd147  : out_data_ref <= 14'h07e2; // 'd2018
      11'd148  : out_data_ref <= 14'h0218; // 'd536
      11'd149  : out_data_ref <= 14'h095a; // 'd2394
      11'd150  : out_data_ref <= 14'h0689; // 'd1673
      11'd151  : out_data_ref <= 14'h08cf; // 'd2255
      11'd152  : out_data_ref <= 14'h069d; // 'd1693
      11'd153  : out_data_ref <= 14'h0248; // 'd584
      11'd154  : out_data_ref <= 14'h09c2; // 'd2498
      11'd155  : out_data_ref <= 14'h014d; // 'd333
      11'd156  : out_data_ref <= 14'h05b1; // 'd1457
      11'd157  : out_data_ref <= 14'h05ed; // 'd1517
      11'd158  : out_data_ref <= 14'h0339; // 'd825
      11'd159  : out_data_ref <= 14'h00ab; // 'd171
      11'd160  : out_data_ref <= 14'h0528; // 'd1320
      11'd161  : out_data_ref <= 14'h08dc; // 'd2268
      11'd162  : out_data_ref <= 14'h02cf; // 'd719
      11'd163  : out_data_ref <= 14'h0414; // 'd1044
      11'd164  : out_data_ref <= 14'h093e; // 'd2366
      11'd165  : out_data_ref <= 14'h0705; // 'd1797
      11'd166  : out_data_ref <= 14'h0894; // 'd2196
      11'd167  : out_data_ref <= 14'h09d9; // 'd2521
      11'd168  : out_data_ref <= 14'h08f9; // 'd2297
      11'd169  : out_data_ref <= 14'h05b9; // 'd1465
      11'd170  : out_data_ref <= 14'h00ae; // 'd174
      11'd171  : out_data_ref <= 14'h0591; // 'd1425
      11'd172  : out_data_ref <= 14'h0318; // 'd792
      11'd173  : out_data_ref <= 14'h061e; // 'd1566
      11'd174  : out_data_ref <= 14'h0a09; // 'd2569
      11'd175  : out_data_ref <= 14'h018a; // 'd394
      11'd176  : out_data_ref <= 14'h09b8; // 'd2488
      11'd177  : out_data_ref <= 14'h03e3; // 'd995
      11'd178  : out_data_ref <= 14'h0998; // 'd2456
      11'd179  : out_data_ref <= 14'h0847; // 'd2119
      11'd180  : out_data_ref <= 14'h0511; // 'd1297
      11'd181  : out_data_ref <= 14'h07ca; // 'd1994
      11'd182  : out_data_ref <= 14'h02b2; // 'd690
      11'd183  : out_data_ref <= 14'h09b9; // 'd2489
      11'd184  : out_data_ref <= 14'h0409; // 'd1033
      11'd185  : out_data_ref <= 14'h06dd; // 'd1757
      11'd186  : out_data_ref <= 14'h011b; // 'd283
      11'd187  : out_data_ref <= 14'h07c9; // 'd1993
      11'd188  : out_data_ref <= 14'h03dc; // 'd988
      11'd189  : out_data_ref <= 14'h0726; // 'd1830
      11'd190  : out_data_ref <= 14'h090c; // 'd2316
      11'd191  : out_data_ref <= 14'h0402; // 'd1026
      11'd192  : out_data_ref <= 14'h0713; // 'd1811
      11'd193  : out_data_ref <= 14'h05b2; // 'd1458
      11'd194  : out_data_ref <= 14'h08e6; // 'd2278
      11'd195  : out_data_ref <= 14'h0201; // 'd513
      11'd196  : out_data_ref <= 14'h04ba; // 'd1210
      11'd197  : out_data_ref <= 14'h04c9; // 'd1225
      11'd198  : out_data_ref <= 14'h048a; // 'd1162
      11'd199  : out_data_ref <= 14'h076f; // 'd1903
      11'd200  : out_data_ref <= 14'h0269; // 'd617
      11'd201  : out_data_ref <= 14'h0572; // 'd1394
      11'd202  : out_data_ref <= 14'h00af; // 'd175
      11'd203  : out_data_ref <= 14'h0315; // 'd789
      11'd204  : out_data_ref <= 14'h0097; // 'd151
      11'd205  : out_data_ref <= 14'h0857; // 'd2135
      11'd206  : out_data_ref <= 14'h098d; // 'd2445
      11'd207  : out_data_ref <= 14'h0134; // 'd308
      11'd208  : out_data_ref <= 14'h00ac; // 'd172
      11'd209  : out_data_ref <= 14'h02d0; // 'd720
      11'd210  : out_data_ref <= 14'h023b; // 'd571
      11'd211  : out_data_ref <= 14'h02a1; // 'd673
      11'd212  : out_data_ref <= 14'h0991; // 'd2449
      11'd213  : out_data_ref <= 14'h01f7; // 'd503
      11'd214  : out_data_ref <= 14'h03cd; // 'd973
      11'd215  : out_data_ref <= 14'h021d; // 'd541
      11'd216  : out_data_ref <= 14'h06ad; // 'd1709
      11'd217  : out_data_ref <= 14'h00fb; // 'd251
      11'd218  : out_data_ref <= 14'h03d5; // 'd981
      11'd219  : out_data_ref <= 14'h0707; // 'd1799
      11'd220  : out_data_ref <= 14'h012e; // 'd302
      11'd221  : out_data_ref <= 14'h0637; // 'd1591
      11'd222  : out_data_ref <= 14'h0786; // 'd1926
      11'd223  : out_data_ref <= 14'h0876; // 'd2166
      11'd224  : out_data_ref <= 14'h00b5; // 'd181
      11'd225  : out_data_ref <= 14'h05ba; // 'd1466
      11'd226  : out_data_ref <= 14'h01ba; // 'd442
      11'd227  : out_data_ref <= 14'h084e; // 'd2126
      11'd228  : out_data_ref <= 14'h067b; // 'd1659
      11'd229  : out_data_ref <= 14'h010f; // 'd271
      11'd230  : out_data_ref <= 14'h070e; // 'd1806
      11'd231  : out_data_ref <= 14'h01f7; // 'd503
      11'd232  : out_data_ref <= 14'h0789; // 'd1929
      11'd233  : out_data_ref <= 14'h04aa; // 'd1194
      11'd234  : out_data_ref <= 14'h0774; // 'd1908
      11'd235  : out_data_ref <= 14'h03a1; // 'd929
      11'd236  : out_data_ref <= 14'h0735; // 'd1845
      11'd237  : out_data_ref <= 14'h0138; // 'd312
      11'd238  : out_data_ref <= 14'h0446; // 'd1094
      11'd239  : out_data_ref <= 14'h02e0; // 'd736
      11'd240  : out_data_ref <= 14'h0942; // 'd2370
      11'd241  : out_data_ref <= 14'h081e; // 'd2078
      11'd242  : out_data_ref <= 14'h0071; // 'd113
      11'd243  : out_data_ref <= 14'h01ad; // 'd429
      11'd244  : out_data_ref <= 14'h0880; // 'd2176
      11'd245  : out_data_ref <= 14'h0159; // 'd345
      11'd246  : out_data_ref <= 14'h0931; // 'd2353
      11'd247  : out_data_ref <= 14'h0756; // 'd1878
      11'd248  : out_data_ref <= 14'h04a1; // 'd1185
      11'd249  : out_data_ref <= 14'h0416; // 'd1046
      11'd250  : out_data_ref <= 14'h03dc; // 'd988
      11'd251  : out_data_ref <= 14'h072a; // 'd1834
      11'd252  : out_data_ref <= 14'h00f2; // 'd242
      11'd253  : out_data_ref <= 14'h02ed; // 'd749
      11'd254  : out_data_ref <= 14'h0664; // 'd1636
      11'd255  : out_data_ref <= 14'h068d; // 'd1677
      11'd256  : out_data_ref <= 14'h04c3; // 'd1219
      11'd257  : out_data_ref <= 14'h0924; // 'd2340
      11'd258  : out_data_ref <= 14'h024e; // 'd590
      11'd259  : out_data_ref <= 14'h0654; // 'd1620
      11'd260  : out_data_ref <= 14'h069e; // 'd1694
      11'd261  : out_data_ref <= 14'h089a; // 'd2202
      11'd262  : out_data_ref <= 14'h06a2; // 'd1698
      11'd263  : out_data_ref <= 14'h05d2; // 'd1490
      11'd264  : out_data_ref <= 14'h01ed; // 'd493
      11'd265  : out_data_ref <= 14'h0273; // 'd627
      11'd266  : out_data_ref <= 14'h0274; // 'd628
      11'd267  : out_data_ref <= 14'h00fb; // 'd251
      11'd268  : out_data_ref <= 14'h072c; // 'd1836
      11'd269  : out_data_ref <= 14'h05f2; // 'd1522
      11'd270  : out_data_ref <= 14'h024e; // 'd590
      11'd271  : out_data_ref <= 14'h0126; // 'd294
      11'd272  : out_data_ref <= 14'h094d; // 'd2381
      11'd273  : out_data_ref <= 14'h0246; // 'd582
      11'd274  : out_data_ref <= 14'h00ce; // 'd206
      11'd275  : out_data_ref <= 14'h0693; // 'd1683
      11'd276  : out_data_ref <= 14'h0983; // 'd2435
      11'd277  : out_data_ref <= 14'h0515; // 'd1301
      11'd278  : out_data_ref <= 14'h06ff; // 'd1791
      11'd279  : out_data_ref <= 14'h055a; // 'd1370
      11'd280  : out_data_ref <= 14'h0259; // 'd601
      11'd281  : out_data_ref <= 14'h0140; // 'd320
      11'd282  : out_data_ref <= 14'h0314; // 'd788
      11'd283  : out_data_ref <= 14'h0706; // 'd1798
      11'd284  : out_data_ref <= 14'h0456; // 'd1110
      11'd285  : out_data_ref <= 14'h0605; // 'd1541
      11'd286  : out_data_ref <= 14'h0296; // 'd662
      11'd287  : out_data_ref <= 14'h06bf; // 'd1727
      11'd288  : out_data_ref <= 14'h04b6; // 'd1206
      11'd289  : out_data_ref <= 14'h075c; // 'd1884
      11'd290  : out_data_ref <= 14'h0564; // 'd1380
      11'd291  : out_data_ref <= 14'h02fb; // 'd763
      11'd292  : out_data_ref <= 14'h03ba; // 'd954
      11'd293  : out_data_ref <= 14'h02fe; // 'd766
      11'd294  : out_data_ref <= 14'h0578; // 'd1400
      11'd295  : out_data_ref <= 14'h0355; // 'd853
      11'd296  : out_data_ref <= 14'h0a00; // 'd2560
      11'd297  : out_data_ref <= 14'h01df; // 'd479
      11'd298  : out_data_ref <= 14'h04ba; // 'd1210
      11'd299  : out_data_ref <= 14'h0052; // 'd82
      11'd300  : out_data_ref <= 14'h0152; // 'd338
      11'd301  : out_data_ref <= 14'h086b; // 'd2155
      11'd302  : out_data_ref <= 14'h0469; // 'd1129
      11'd303  : out_data_ref <= 14'h07f3; // 'd2035
      11'd304  : out_data_ref <= 14'h038c; // 'd908
      11'd305  : out_data_ref <= 14'h0102; // 'd258
      11'd306  : out_data_ref <= 14'h00ec; // 'd236
      11'd307  : out_data_ref <= 14'h06f9; // 'd1785
      11'd308  : out_data_ref <= 14'h04fd; // 'd1277
      11'd309  : out_data_ref <= 14'h0991; // 'd2449
      11'd310  : out_data_ref <= 14'h0470; // 'd1136
      11'd311  : out_data_ref <= 14'h032d; // 'd813
      11'd312  : out_data_ref <= 14'h083d; // 'd2109
      11'd313  : out_data_ref <= 14'h0099; // 'd153
      11'd314  : out_data_ref <= 14'h01c4; // 'd452
      11'd315  : out_data_ref <= 14'h0303; // 'd771
      11'd316  : out_data_ref <= 14'h08a3; // 'd2211
      11'd317  : out_data_ref <= 14'h01cd; // 'd461
      11'd318  : out_data_ref <= 14'h057f; // 'd1407
      11'd319  : out_data_ref <= 14'h0996; // 'd2454
      11'd320  : out_data_ref <= 14'h04fc; // 'd1276
      11'd321  : out_data_ref <= 14'h049b; // 'd1179
      11'd322  : out_data_ref <= 14'h0899; // 'd2201
      11'd323  : out_data_ref <= 14'h04d4; // 'd1236
      11'd324  : out_data_ref <= 14'h0a02; // 'd2562
      11'd325  : out_data_ref <= 14'h06e5; // 'd1765
      11'd326  : out_data_ref <= 14'h08ff; // 'd2303
      11'd327  : out_data_ref <= 14'h07cb; // 'd1995
      11'd328  : out_data_ref <= 14'h0803; // 'd2051
      11'd329  : out_data_ref <= 14'h0392; // 'd914
      11'd330  : out_data_ref <= 14'h0186; // 'd390
      11'd331  : out_data_ref <= 14'h0285; // 'd645
      11'd332  : out_data_ref <= 14'h07de; // 'd2014
      11'd333  : out_data_ref <= 14'h00bc; // 'd188
      11'd334  : out_data_ref <= 14'h07eb; // 'd2027
      11'd335  : out_data_ref <= 14'h063f; // 'd1599
      11'd336  : out_data_ref <= 14'h091e; // 'd2334
      11'd337  : out_data_ref <= 14'h009a; // 'd154
      11'd338  : out_data_ref <= 14'h07f5; // 'd2037
      11'd339  : out_data_ref <= 14'h050e; // 'd1294
      11'd340  : out_data_ref <= 14'h0799; // 'd1945
      11'd341  : out_data_ref <= 14'h04e8; // 'd1256
      11'd342  : out_data_ref <= 14'h0a0d; // 'd2573
      11'd343  : out_data_ref <= 14'h04a7; // 'd1191
      11'd344  : out_data_ref <= 14'h096f; // 'd2415
      11'd345  : out_data_ref <= 14'h090e; // 'd2318
      11'd346  : out_data_ref <= 14'h068a; // 'd1674
      11'd347  : out_data_ref <= 14'h079c; // 'd1948
      11'd348  : out_data_ref <= 14'h08cd; // 'd2253
      11'd349  : out_data_ref <= 14'h0293; // 'd659
      11'd350  : out_data_ref <= 14'h04dd; // 'd1245
      11'd351  : out_data_ref <= 14'h0805; // 'd2053
      11'd352  : out_data_ref <= 14'h0402; // 'd1026
      11'd353  : out_data_ref <= 14'h016e; // 'd366
      11'd354  : out_data_ref <= 14'h0454; // 'd1108
      11'd355  : out_data_ref <= 14'h06cc; // 'd1740
      11'd356  : out_data_ref <= 14'h0675; // 'd1653
      11'd357  : out_data_ref <= 14'h03be; // 'd958
      11'd358  : out_data_ref <= 14'h0889; // 'd2185
      11'd359  : out_data_ref <= 14'h0843; // 'd2115
      11'd360  : out_data_ref <= 14'h0762; // 'd1890
      11'd361  : out_data_ref <= 14'h03ad; // 'd941
      11'd362  : out_data_ref <= 14'h055c; // 'd1372
      11'd363  : out_data_ref <= 14'h0a1e; // 'd2590
      11'd364  : out_data_ref <= 14'h075f; // 'd1887
      11'd365  : out_data_ref <= 14'h0495; // 'd1173
      11'd366  : out_data_ref <= 14'h063b; // 'd1595
      11'd367  : out_data_ref <= 14'h022a; // 'd554
      11'd368  : out_data_ref <= 14'h050a; // 'd1290
      11'd369  : out_data_ref <= 14'h06d7; // 'd1751
      11'd370  : out_data_ref <= 14'h0248; // 'd584
      11'd371  : out_data_ref <= 14'h01c3; // 'd451
      11'd372  : out_data_ref <= 14'h05a9; // 'd1449
      11'd373  : out_data_ref <= 14'h0599; // 'd1433
      11'd374  : out_data_ref <= 14'h0028; // 'd40
      11'd375  : out_data_ref <= 14'h00cb; // 'd203
      11'd376  : out_data_ref <= 14'h0237; // 'd567
      11'd377  : out_data_ref <= 14'h04ca; // 'd1226
      11'd378  : out_data_ref <= 14'h007d; // 'd125
      11'd379  : out_data_ref <= 14'h05d2; // 'd1490
      11'd380  : out_data_ref <= 14'h0005; // 'd5
      11'd381  : out_data_ref <= 14'h0415; // 'd1045
      11'd382  : out_data_ref <= 14'h016c; // 'd364
      11'd383  : out_data_ref <= 14'h09a4; // 'd2468
      11'd384  : out_data_ref <= 14'h06d0; // 'd1744
      11'd385  : out_data_ref <= 14'h0999; // 'd2457
      11'd386  : out_data_ref <= 14'h08d8; // 'd2264
      11'd387  : out_data_ref <= 14'h06a8; // 'd1704
      11'd388  : out_data_ref <= 14'h03c0; // 'd960
      11'd389  : out_data_ref <= 14'h0181; // 'd385
      11'd390  : out_data_ref <= 14'h0142; // 'd322
      11'd391  : out_data_ref <= 14'h096f; // 'd2415
      11'd392  : out_data_ref <= 14'h069a; // 'd1690
      11'd393  : out_data_ref <= 14'h015d; // 'd349
      11'd394  : out_data_ref <= 14'h0594; // 'd1428
      11'd395  : out_data_ref <= 14'h090d; // 'd2317
      11'd396  : out_data_ref <= 14'h063a; // 'd1594
      11'd397  : out_data_ref <= 14'h09fb; // 'd2555
      11'd398  : out_data_ref <= 14'h00a2; // 'd162
      11'd399  : out_data_ref <= 14'h0523; // 'd1315
      11'd400  : out_data_ref <= 14'h05eb; // 'd1515
      11'd401  : out_data_ref <= 14'h041b; // 'd1051
      11'd402  : out_data_ref <= 14'h0955; // 'd2389
      11'd403  : out_data_ref <= 14'h006f; // 'd111
      11'd404  : out_data_ref <= 14'h04eb; // 'd1259
      11'd405  : out_data_ref <= 14'h05de; // 'd1502
      11'd406  : out_data_ref <= 14'h057b; // 'd1403
      11'd407  : out_data_ref <= 14'h032a; // 'd810
      11'd408  : out_data_ref <= 14'h073f; // 'd1855
      11'd409  : out_data_ref <= 14'h0943; // 'd2371
      11'd410  : out_data_ref <= 14'h05eb; // 'd1515
      11'd411  : out_data_ref <= 14'h08c1; // 'd2241
      11'd412  : out_data_ref <= 14'h011d; // 'd285
      11'd413  : out_data_ref <= 14'h0658; // 'd1624
      11'd414  : out_data_ref <= 14'h03d3; // 'd979
      11'd415  : out_data_ref <= 14'h01f6; // 'd502
      11'd416  : out_data_ref <= 14'h0671; // 'd1649
      11'd417  : out_data_ref <= 14'h0089; // 'd137
      11'd418  : out_data_ref <= 14'h0117; // 'd279
      11'd419  : out_data_ref <= 14'h04a6; // 'd1190
      11'd420  : out_data_ref <= 14'h07e2; // 'd2018
      11'd421  : out_data_ref <= 14'h032a; // 'd810
      11'd422  : out_data_ref <= 14'h06b1; // 'd1713
      11'd423  : out_data_ref <= 14'h0825; // 'd2085
      11'd424  : out_data_ref <= 14'h0086; // 'd134
      11'd425  : out_data_ref <= 14'h012a; // 'd298
      11'd426  : out_data_ref <= 14'h05d7; // 'd1495
      11'd427  : out_data_ref <= 14'h0680; // 'd1664
      11'd428  : out_data_ref <= 14'h05c2; // 'd1474
      11'd429  : out_data_ref <= 14'h01df; // 'd479
      11'd430  : out_data_ref <= 14'h031a; // 'd794
      11'd431  : out_data_ref <= 14'h09c6; // 'd2502
      11'd432  : out_data_ref <= 14'h03cb; // 'd971
      11'd433  : out_data_ref <= 14'h0408; // 'd1032
      11'd434  : out_data_ref <= 14'h0007; // 'd7
      11'd435  : out_data_ref <= 14'h06be; // 'd1726
      11'd436  : out_data_ref <= 14'h07ea; // 'd2026
      11'd437  : out_data_ref <= 14'h095b; // 'd2395
      11'd438  : out_data_ref <= 14'h09d6; // 'd2518
      11'd439  : out_data_ref <= 14'h09bf; // 'd2495
      11'd440  : out_data_ref <= 14'h097c; // 'd2428
      11'd441  : out_data_ref <= 14'h0416; // 'd1046
      11'd442  : out_data_ref <= 14'h04cc; // 'd1228
      11'd443  : out_data_ref <= 14'h08c4; // 'd2244
      11'd444  : out_data_ref <= 14'h064b; // 'd1611
      11'd445  : out_data_ref <= 14'h059d; // 'd1437
      11'd446  : out_data_ref <= 14'h0278; // 'd632
      11'd447  : out_data_ref <= 14'h00e8; // 'd232
      11'd448  : out_data_ref <= 14'h0834; // 'd2100
      11'd449  : out_data_ref <= 14'h03de; // 'd990
      11'd450  : out_data_ref <= 14'h0233; // 'd563
      11'd451  : out_data_ref <= 14'h09db; // 'd2523
      11'd452  : out_data_ref <= 14'h02c5; // 'd709
      11'd453  : out_data_ref <= 14'h08d6; // 'd2262
      11'd454  : out_data_ref <= 14'h050a; // 'd1290
      11'd455  : out_data_ref <= 14'h0636; // 'd1590
      11'd456  : out_data_ref <= 14'h023b; // 'd571
      11'd457  : out_data_ref <= 14'h009b; // 'd155
      11'd458  : out_data_ref <= 14'h004f; // 'd79
      11'd459  : out_data_ref <= 14'h0408; // 'd1032
      11'd460  : out_data_ref <= 14'h014a; // 'd330
      11'd461  : out_data_ref <= 14'h03ea; // 'd1002
      11'd462  : out_data_ref <= 14'h08e4; // 'd2276
      11'd463  : out_data_ref <= 14'h0398; // 'd920
      11'd464  : out_data_ref <= 14'h0716; // 'd1814
      11'd465  : out_data_ref <= 14'h0212; // 'd530
      11'd466  : out_data_ref <= 14'h0563; // 'd1379
      11'd467  : out_data_ref <= 14'h07d2; // 'd2002
      11'd468  : out_data_ref <= 14'h01e3; // 'd483
      11'd469  : out_data_ref <= 14'h04b3; // 'd1203
      11'd470  : out_data_ref <= 14'h021a; // 'd538
      11'd471  : out_data_ref <= 14'h0423; // 'd1059
      11'd472  : out_data_ref <= 14'h01f3; // 'd499
      11'd473  : out_data_ref <= 14'h0230; // 'd560
      11'd474  : out_data_ref <= 14'h045a; // 'd1114
      11'd475  : out_data_ref <= 14'h0025; // 'd37
      11'd476  : out_data_ref <= 14'h026f; // 'd623
      11'd477  : out_data_ref <= 14'h0004; // 'd4
      11'd478  : out_data_ref <= 14'h00f9; // 'd249
      11'd479  : out_data_ref <= 14'h00e7; // 'd231
      11'd480  : out_data_ref <= 14'h0a3b; // 'd2619
      11'd481  : out_data_ref <= 14'h0426; // 'd1062
      11'd482  : out_data_ref <= 14'h01a5; // 'd421
      11'd483  : out_data_ref <= 14'h02a0; // 'd672
      11'd484  : out_data_ref <= 14'h060d; // 'd1549
      11'd485  : out_data_ref <= 14'h0707; // 'd1799
      11'd486  : out_data_ref <= 14'h010a; // 'd266
      11'd487  : out_data_ref <= 14'h03e2; // 'd994
      11'd488  : out_data_ref <= 14'h0583; // 'd1411
      11'd489  : out_data_ref <= 14'h031c; // 'd796
      11'd490  : out_data_ref <= 14'h08e1; // 'd2273
      11'd491  : out_data_ref <= 14'h0a35; // 'd2613
      11'd492  : out_data_ref <= 14'h071e; // 'd1822
      11'd493  : out_data_ref <= 14'h06c2; // 'd1730
      11'd494  : out_data_ref <= 14'h0688; // 'd1672
      11'd495  : out_data_ref <= 14'h0134; // 'd308
      11'd496  : out_data_ref <= 14'h0461; // 'd1121
      11'd497  : out_data_ref <= 14'h06b5; // 'd1717
      11'd498  : out_data_ref <= 14'h0729; // 'd1833
      11'd499  : out_data_ref <= 14'h06e0; // 'd1760
      11'd500  : out_data_ref <= 14'h0737; // 'd1847
      11'd501  : out_data_ref <= 14'h07fd; // 'd2045
      11'd502  : out_data_ref <= 14'h000f; // 'd15
      11'd503  : out_data_ref <= 14'h04d1; // 'd1233
      11'd504  : out_data_ref <= 14'h0248; // 'd584
      11'd505  : out_data_ref <= 14'h0635; // 'd1589
      11'd506  : out_data_ref <= 14'h0988; // 'd2440
      11'd507  : out_data_ref <= 14'h075f; // 'd1887
      11'd508  : out_data_ref <= 14'h0310; // 'd784
      11'd509  : out_data_ref <= 14'h086d; // 'd2157
      11'd510  : out_data_ref <= 14'h0828; // 'd2088
      11'd511  : out_data_ref <= 14'h022c; // 'd556
      11'd512  : out_data_ref <= 14'h0283; // 'd643
      11'd513  : out_data_ref <= 14'h0a24; // 'd2596
      11'd514  : out_data_ref <= 14'h046a; // 'd1130
      11'd515  : out_data_ref <= 14'h09fd; // 'd2557
      11'd516  : out_data_ref <= 14'h05fa; // 'd1530
      11'd517  : out_data_ref <= 14'h082b; // 'd2091
      11'd518  : out_data_ref <= 14'h02d7; // 'd727
      11'd519  : out_data_ref <= 14'h06f4; // 'd1780
      11'd520  : out_data_ref <= 14'h0a30; // 'd2608
      11'd521  : out_data_ref <= 14'h0693; // 'd1683
      11'd522  : out_data_ref <= 14'h02fb; // 'd763
      11'd523  : out_data_ref <= 14'h09bf; // 'd2495
      11'd524  : out_data_ref <= 14'h04cf; // 'd1231
      11'd525  : out_data_ref <= 14'h021f; // 'd543
      11'd526  : out_data_ref <= 14'h04be; // 'd1214
      11'd527  : out_data_ref <= 14'h039d; // 'd925
      11'd528  : out_data_ref <= 14'h05fa; // 'd1530
      11'd529  : out_data_ref <= 14'h05a6; // 'd1446
      11'd530  : out_data_ref <= 14'h0128; // 'd296
      11'd531  : out_data_ref <= 14'h0961; // 'd2401
      11'd532  : out_data_ref <= 14'h01ce; // 'd462
      11'd533  : out_data_ref <= 14'h05b3; // 'd1459
      11'd534  : out_data_ref <= 14'h03b4; // 'd948
      11'd535  : out_data_ref <= 14'h097a; // 'd2426
      11'd536  : out_data_ref <= 14'h065c; // 'd1628
      11'd537  : out_data_ref <= 14'h0479; // 'd1145
      11'd538  : out_data_ref <= 14'h0574; // 'd1396
      11'd539  : out_data_ref <= 14'h0a27; // 'd2599
      11'd540  : out_data_ref <= 14'h04cf; // 'd1231
      11'd541  : out_data_ref <= 14'h038e; // 'd910
      11'd542  : out_data_ref <= 14'h0520; // 'd1312
      11'd543  : out_data_ref <= 14'h01b9; // 'd441
      11'd544  : out_data_ref <= 14'h0a03; // 'd2563
      11'd545  : out_data_ref <= 14'h0988; // 'd2440
      11'd546  : out_data_ref <= 14'h0227; // 'd551
      11'd547  : out_data_ref <= 14'h056d; // 'd1389
      11'd548  : out_data_ref <= 14'h0230; // 'd560
      11'd549  : out_data_ref <= 14'h03f6; // 'd1014
      11'd550  : out_data_ref <= 14'h08a2; // 'd2210
      11'd551  : out_data_ref <= 14'h0277; // 'd631
      11'd552  : out_data_ref <= 14'h08c8; // 'd2248
      11'd553  : out_data_ref <= 14'h003f; // 'd63
      11'd554  : out_data_ref <= 14'h0951; // 'd2385
      11'd555  : out_data_ref <= 14'h04d0; // 'd1232
      11'd556  : out_data_ref <= 14'h091a; // 'd2330
      11'd557  : out_data_ref <= 14'h0985; // 'd2437
      11'd558  : out_data_ref <= 14'h032f; // 'd815
      11'd559  : out_data_ref <= 14'h044c; // 'd1100
      11'd560  : out_data_ref <= 14'h075d; // 'd1885
      11'd561  : out_data_ref <= 14'h05a6; // 'd1446
      11'd562  : out_data_ref <= 14'h0286; // 'd646
      11'd563  : out_data_ref <= 14'h040f; // 'd1039
      11'd564  : out_data_ref <= 14'h013c; // 'd316
      11'd565  : out_data_ref <= 14'h0a1f; // 'd2591
      11'd566  : out_data_ref <= 14'h08d9; // 'd2265
      11'd567  : out_data_ref <= 14'h07a1; // 'd1953
      11'd568  : out_data_ref <= 14'h03ca; // 'd970
      11'd569  : out_data_ref <= 14'h0368; // 'd872
      11'd570  : out_data_ref <= 14'h06e8; // 'd1768
      11'd571  : out_data_ref <= 14'h03cb; // 'd971
      11'd572  : out_data_ref <= 14'h029a; // 'd666
      11'd573  : out_data_ref <= 14'h08db; // 'd2267
      11'd574  : out_data_ref <= 14'h059e; // 'd1438
      11'd575  : out_data_ref <= 14'h0767; // 'd1895
      11'd576  : out_data_ref <= 14'h02c2; // 'd706
      11'd577  : out_data_ref <= 14'h07f1; // 'd2033
      11'd578  : out_data_ref <= 14'h01cc; // 'd460
      11'd579  : out_data_ref <= 14'h0286; // 'd646
      11'd580  : out_data_ref <= 14'h0068; // 'd104
      11'd581  : out_data_ref <= 14'h079b; // 'd1947
      11'd582  : out_data_ref <= 14'h010d; // 'd269
      11'd583  : out_data_ref <= 14'h051a; // 'd1306
      11'd584  : out_data_ref <= 14'h01f5; // 'd501
      11'd585  : out_data_ref <= 14'h002b; // 'd43
      11'd586  : out_data_ref <= 14'h0738; // 'd1848
      11'd587  : out_data_ref <= 14'h0399; // 'd921
      11'd588  : out_data_ref <= 14'h0562; // 'd1378
      11'd589  : out_data_ref <= 14'h03d6; // 'd982
      11'd590  : out_data_ref <= 14'h0232; // 'd562
      11'd591  : out_data_ref <= 14'h0811; // 'd2065
      11'd592  : out_data_ref <= 14'h003a; // 'd58
      11'd593  : out_data_ref <= 14'h0649; // 'd1609
      11'd594  : out_data_ref <= 14'h016d; // 'd365
      11'd595  : out_data_ref <= 14'h0079; // 'd121
      11'd596  : out_data_ref <= 14'h091e; // 'd2334
      11'd597  : out_data_ref <= 14'h045d; // 'd1117
      11'd598  : out_data_ref <= 14'h07f6; // 'd2038
      11'd599  : out_data_ref <= 14'h06dc; // 'd1756
      11'd600  : out_data_ref <= 14'h001d; // 'd29
      11'd601  : out_data_ref <= 14'h03a8; // 'd936
      11'd602  : out_data_ref <= 14'h053f; // 'd1343
      11'd603  : out_data_ref <= 14'h044a; // 'd1098
      11'd604  : out_data_ref <= 14'h06b3; // 'd1715
      11'd605  : out_data_ref <= 14'h02b6; // 'd694
      11'd606  : out_data_ref <= 14'h03eb; // 'd1003
      11'd607  : out_data_ref <= 14'h00cf; // 'd207
      11'd608  : out_data_ref <= 14'h06f1; // 'd1777
      11'd609  : out_data_ref <= 14'h0138; // 'd312
      11'd610  : out_data_ref <= 14'h012a; // 'd298
      11'd611  : out_data_ref <= 14'h0275; // 'd629
      11'd612  : out_data_ref <= 14'h0259; // 'd601
      11'd613  : out_data_ref <= 14'h0699; // 'd1689
      11'd614  : out_data_ref <= 14'h08c8; // 'd2248
      11'd615  : out_data_ref <= 14'h08ef; // 'd2287
      11'd616  : out_data_ref <= 14'h0255; // 'd597
      11'd617  : out_data_ref <= 14'h0032; // 'd50
      11'd618  : out_data_ref <= 14'h06bc; // 'd1724
      11'd619  : out_data_ref <= 14'h0242; // 'd578
      11'd620  : out_data_ref <= 14'h0803; // 'd2051
      11'd621  : out_data_ref <= 14'h0542; // 'd1346
      11'd622  : out_data_ref <= 14'h015b; // 'd347
      11'd623  : out_data_ref <= 14'h0980; // 'd2432
      11'd624  : out_data_ref <= 14'h0988; // 'd2440
      11'd625  : out_data_ref <= 14'h0628; // 'd1576
      11'd626  : out_data_ref <= 14'h07fc; // 'd2044
      11'd627  : out_data_ref <= 14'h0988; // 'd2440
      11'd628  : out_data_ref <= 14'h067a; // 'd1658
      11'd629  : out_data_ref <= 14'h0a3d; // 'd2621
      11'd630  : out_data_ref <= 14'h00a1; // 'd161
      11'd631  : out_data_ref <= 14'h097e; // 'd2430
      11'd632  : out_data_ref <= 14'h00a8; // 'd168
      11'd633  : out_data_ref <= 14'h09a3; // 'd2467
      11'd634  : out_data_ref <= 14'h05a0; // 'd1440
      11'd635  : out_data_ref <= 14'h0738; // 'd1848
      11'd636  : out_data_ref <= 14'h0412; // 'd1042
      11'd637  : out_data_ref <= 14'h09c9; // 'd2505
      11'd638  : out_data_ref <= 14'h0987; // 'd2439
      11'd639  : out_data_ref <= 14'h0070; // 'd112
      11'd640  : out_data_ref <= 14'h0369; // 'd873
      11'd641  : out_data_ref <= 14'h0587; // 'd1415
      11'd642  : out_data_ref <= 14'h07a6; // 'd1958
      11'd643  : out_data_ref <= 14'h0233; // 'd563
      11'd644  : out_data_ref <= 14'h0731; // 'd1841
      11'd645  : out_data_ref <= 14'h0116; // 'd278
      11'd646  : out_data_ref <= 14'h03aa; // 'd938
      11'd647  : out_data_ref <= 14'h00f6; // 'd246
      11'd648  : out_data_ref <= 14'h040d; // 'd1037
      11'd649  : out_data_ref <= 14'h0335; // 'd821
      11'd650  : out_data_ref <= 14'h0936; // 'd2358
      11'd651  : out_data_ref <= 14'h0950; // 'd2384
      11'd652  : out_data_ref <= 14'h0736; // 'd1846
      11'd653  : out_data_ref <= 14'h001f; // 'd31
      11'd654  : out_data_ref <= 14'h02e5; // 'd741
      11'd655  : out_data_ref <= 14'h08d1; // 'd2257
      11'd656  : out_data_ref <= 14'h07be; // 'd1982
      11'd657  : out_data_ref <= 14'h0240; // 'd576
      11'd658  : out_data_ref <= 14'h06a3; // 'd1699
      11'd659  : out_data_ref <= 14'h07e2; // 'd2018
      11'd660  : out_data_ref <= 14'h010c; // 'd268
      11'd661  : out_data_ref <= 14'h0271; // 'd625
      11'd662  : out_data_ref <= 14'h0167; // 'd359
      11'd663  : out_data_ref <= 14'h040c; // 'd1036
      11'd664  : out_data_ref <= 14'h06f0; // 'd1776
      11'd665  : out_data_ref <= 14'h00b5; // 'd181
      11'd666  : out_data_ref <= 14'h07a1; // 'd1953
      11'd667  : out_data_ref <= 14'h017d; // 'd381
      11'd668  : out_data_ref <= 14'h0262; // 'd610
      11'd669  : out_data_ref <= 14'h090e; // 'd2318
      11'd670  : out_data_ref <= 14'h0522; // 'd1314
      11'd671  : out_data_ref <= 14'h05cb; // 'd1483
      11'd672  : out_data_ref <= 14'h03cc; // 'd972
      11'd673  : out_data_ref <= 14'h02a3; // 'd675
      11'd674  : out_data_ref <= 14'h0166; // 'd358
      11'd675  : out_data_ref <= 14'h007d; // 'd125
      11'd676  : out_data_ref <= 14'h01de; // 'd478
      11'd677  : out_data_ref <= 14'h0250; // 'd592
      11'd678  : out_data_ref <= 14'h04df; // 'd1247
      11'd679  : out_data_ref <= 14'h033b; // 'd827
      11'd680  : out_data_ref <= 14'h085d; // 'd2141
      11'd681  : out_data_ref <= 14'h022a; // 'd554
      11'd682  : out_data_ref <= 14'h0750; // 'd1872
      11'd683  : out_data_ref <= 14'h0178; // 'd376
      11'd684  : out_data_ref <= 14'h03ee; // 'd1006
      11'd685  : out_data_ref <= 14'h0073; // 'd115
      11'd686  : out_data_ref <= 14'h0642; // 'd1602
      11'd687  : out_data_ref <= 14'h03f4; // 'd1012
      11'd688  : out_data_ref <= 14'h01b9; // 'd441
      11'd689  : out_data_ref <= 14'h0708; // 'd1800
      11'd690  : out_data_ref <= 14'h0843; // 'd2115
      11'd691  : out_data_ref <= 14'h06d5; // 'd1749
      11'd692  : out_data_ref <= 14'h014d; // 'd333
      11'd693  : out_data_ref <= 14'h0564; // 'd1380
      11'd694  : out_data_ref <= 14'h01bc; // 'd444
      11'd695  : out_data_ref <= 14'h00e2; // 'd226
      11'd696  : out_data_ref <= 14'h0750; // 'd1872
      11'd697  : out_data_ref <= 14'h07f7; // 'd2039
      11'd698  : out_data_ref <= 14'h0453; // 'd1107
      11'd699  : out_data_ref <= 14'h05da; // 'd1498
      11'd700  : out_data_ref <= 14'h0868; // 'd2152
      11'd701  : out_data_ref <= 14'h000d; // 'd13
      11'd702  : out_data_ref <= 14'h0a40; // 'd2624
      11'd703  : out_data_ref <= 14'h0963; // 'd2403
      11'd704  : out_data_ref <= 14'h0801; // 'd2049
      11'd705  : out_data_ref <= 14'h07e1; // 'd2017
      11'd706  : out_data_ref <= 14'h02d9; // 'd729
      11'd707  : out_data_ref <= 14'h0406; // 'd1030
      11'd708  : out_data_ref <= 14'h0328; // 'd808
      11'd709  : out_data_ref <= 14'h01af; // 'd431
      11'd710  : out_data_ref <= 14'h04b6; // 'd1206
      11'd711  : out_data_ref <= 14'h03ea; // 'd1002
      11'd712  : out_data_ref <= 14'h02fa; // 'd762
      11'd713  : out_data_ref <= 14'h04dc; // 'd1244
      11'd714  : out_data_ref <= 14'h02fb; // 'd763
      11'd715  : out_data_ref <= 14'h040c; // 'd1036
      11'd716  : out_data_ref <= 14'h068a; // 'd1674
      11'd717  : out_data_ref <= 14'h086c; // 'd2156
      11'd718  : out_data_ref <= 14'h043b; // 'd1083
      11'd719  : out_data_ref <= 14'h0816; // 'd2070
      11'd720  : out_data_ref <= 14'h0270; // 'd624
      11'd721  : out_data_ref <= 14'h0224; // 'd548
      11'd722  : out_data_ref <= 14'h0809; // 'd2057
      11'd723  : out_data_ref <= 14'h09d5; // 'd2517
      11'd724  : out_data_ref <= 14'h012c; // 'd300
      11'd725  : out_data_ref <= 14'h08dc; // 'd2268
      11'd726  : out_data_ref <= 14'h02f4; // 'd756
      11'd727  : out_data_ref <= 14'h06b0; // 'd1712
      11'd728  : out_data_ref <= 14'h022f; // 'd559
      11'd729  : out_data_ref <= 14'h035a; // 'd858
      11'd730  : out_data_ref <= 14'h0473; // 'd1139
      11'd731  : out_data_ref <= 14'h0136; // 'd310
      11'd732  : out_data_ref <= 14'h09c9; // 'd2505
      11'd733  : out_data_ref <= 14'h08cf; // 'd2255
      11'd734  : out_data_ref <= 14'h0684; // 'd1668
      11'd735  : out_data_ref <= 14'h08df; // 'd2271
      11'd736  : out_data_ref <= 14'h078a; // 'd1930
      11'd737  : out_data_ref <= 14'h078c; // 'd1932
      11'd738  : out_data_ref <= 14'h0682; // 'd1666
      11'd739  : out_data_ref <= 14'h0253; // 'd595
      11'd740  : out_data_ref <= 14'h04f2; // 'd1266
      11'd741  : out_data_ref <= 14'h06ff; // 'd1791
      11'd742  : out_data_ref <= 14'h006b; // 'd107
      11'd743  : out_data_ref <= 14'h0453; // 'd1107
      11'd744  : out_data_ref <= 14'h0109; // 'd265
      11'd745  : out_data_ref <= 14'h037c; // 'd892
      11'd746  : out_data_ref <= 14'h0838; // 'd2104
      11'd747  : out_data_ref <= 14'h03c8; // 'd968
      11'd748  : out_data_ref <= 14'h0564; // 'd1380
      11'd749  : out_data_ref <= 14'h06c7; // 'd1735
      11'd750  : out_data_ref <= 14'h0581; // 'd1409
      11'd751  : out_data_ref <= 14'h036c; // 'd876
      11'd752  : out_data_ref <= 14'h0034; // 'd52
      11'd753  : out_data_ref <= 14'h07a8; // 'd1960
      11'd754  : out_data_ref <= 14'h055a; // 'd1370
      11'd755  : out_data_ref <= 14'h0271; // 'd625
      11'd756  : out_data_ref <= 14'h038b; // 'd907
      11'd757  : out_data_ref <= 14'h09b2; // 'd2482
      11'd758  : out_data_ref <= 14'h037a; // 'd890
      11'd759  : out_data_ref <= 14'h0991; // 'd2449
      11'd760  : out_data_ref <= 14'h0712; // 'd1810
      11'd761  : out_data_ref <= 14'h0890; // 'd2192
      11'd762  : out_data_ref <= 14'h01cb; // 'd459
      11'd763  : out_data_ref <= 14'h086b; // 'd2155
      11'd764  : out_data_ref <= 14'h066f; // 'd1647
      11'd765  : out_data_ref <= 14'h06bf; // 'd1727
      11'd766  : out_data_ref <= 14'h01bc; // 'd444
      11'd767  : out_data_ref <= 14'h010d; // 'd269
      11'd768  : out_data_ref <= 14'h082d; // 'd2093
      11'd769  : out_data_ref <= 14'h094a; // 'd2378
      11'd770  : out_data_ref <= 14'h06f2; // 'd1778
      11'd771  : out_data_ref <= 14'h067a; // 'd1658
      11'd772  : out_data_ref <= 14'h05c4; // 'd1476
      11'd773  : out_data_ref <= 14'h03c4; // 'd964
      11'd774  : out_data_ref <= 14'h0598; // 'd1432
      11'd775  : out_data_ref <= 14'h0402; // 'd1026
      11'd776  : out_data_ref <= 14'h01a8; // 'd424
      11'd777  : out_data_ref <= 14'h0152; // 'd338
      11'd778  : out_data_ref <= 14'h068e; // 'd1678
      11'd779  : out_data_ref <= 14'h09d1; // 'd2513
      11'd780  : out_data_ref <= 14'h081e; // 'd2078
      11'd781  : out_data_ref <= 14'h06fd; // 'd1789
      11'd782  : out_data_ref <= 14'h0861; // 'd2145
      11'd783  : out_data_ref <= 14'h072c; // 'd1836
      11'd784  : out_data_ref <= 14'h0842; // 'd2114
      11'd785  : out_data_ref <= 14'h085c; // 'd2140
      11'd786  : out_data_ref <= 14'h0429; // 'd1065
      11'd787  : out_data_ref <= 14'h0314; // 'd788
      11'd788  : out_data_ref <= 14'h01bd; // 'd445
      11'd789  : out_data_ref <= 14'h09e5; // 'd2533
      11'd790  : out_data_ref <= 14'h06fb; // 'd1787
      11'd791  : out_data_ref <= 14'h0929; // 'd2345
      11'd792  : out_data_ref <= 14'h07ce; // 'd1998
      11'd793  : out_data_ref <= 14'h06b4; // 'd1716
      11'd794  : out_data_ref <= 14'h0350; // 'd848
      11'd795  : out_data_ref <= 14'h0991; // 'd2449
      11'd796  : out_data_ref <= 14'h05f8; // 'd1528
      11'd797  : out_data_ref <= 14'h02ed; // 'd749
      11'd798  : out_data_ref <= 14'h04d3; // 'd1235
      11'd799  : out_data_ref <= 14'h0358; // 'd856
      11'd800  : out_data_ref <= 14'h010e; // 'd270
      11'd801  : out_data_ref <= 14'h0742; // 'd1858
      11'd802  : out_data_ref <= 14'h05b5; // 'd1461
      11'd803  : out_data_ref <= 14'h00da; // 'd218
      11'd804  : out_data_ref <= 14'h039e; // 'd926
      11'd805  : out_data_ref <= 14'h051f; // 'd1311
      11'd806  : out_data_ref <= 14'h0055; // 'd85
      11'd807  : out_data_ref <= 14'h0571; // 'd1393
      11'd808  : out_data_ref <= 14'h057d; // 'd1405
      11'd809  : out_data_ref <= 14'h0028; // 'd40
      11'd810  : out_data_ref <= 14'h0a02; // 'd2562
      11'd811  : out_data_ref <= 14'h0066; // 'd102
      11'd812  : out_data_ref <= 14'h073c; // 'd1852
      11'd813  : out_data_ref <= 14'h0788; // 'd1928
      11'd814  : out_data_ref <= 14'h016a; // 'd362
      11'd815  : out_data_ref <= 14'h08e4; // 'd2276
      11'd816  : out_data_ref <= 14'h01a4; // 'd420
      11'd817  : out_data_ref <= 14'h089e; // 'd2206
      11'd818  : out_data_ref <= 14'h08bb; // 'd2235
      11'd819  : out_data_ref <= 14'h0597; // 'd1431
      11'd820  : out_data_ref <= 14'h026d; // 'd621
      11'd821  : out_data_ref <= 14'h00a4; // 'd164
      11'd822  : out_data_ref <= 14'h0602; // 'd1538
      11'd823  : out_data_ref <= 14'h07b7; // 'd1975
      11'd824  : out_data_ref <= 14'h06ce; // 'd1742
      11'd825  : out_data_ref <= 14'h0a01; // 'd2561
      11'd826  : out_data_ref <= 14'h071d; // 'd1821
      11'd827  : out_data_ref <= 14'h09be; // 'd2494
      11'd828  : out_data_ref <= 14'h0018; // 'd24
      11'd829  : out_data_ref <= 14'h0119; // 'd281
      11'd830  : out_data_ref <= 14'h0390; // 'd912
      11'd831  : out_data_ref <= 14'h04c5; // 'd1221
      11'd832  : out_data_ref <= 14'h0112; // 'd274
      11'd833  : out_data_ref <= 14'h005d; // 'd93
      11'd834  : out_data_ref <= 14'h08ec; // 'd2284
      11'd835  : out_data_ref <= 14'h00ad; // 'd173
      11'd836  : out_data_ref <= 14'h02b5; // 'd693
      11'd837  : out_data_ref <= 14'h08b0; // 'd2224
      11'd838  : out_data_ref <= 14'h0317; // 'd791
      11'd839  : out_data_ref <= 14'h0088; // 'd136
      11'd840  : out_data_ref <= 14'h09eb; // 'd2539
      11'd841  : out_data_ref <= 14'h03a8; // 'd936
      11'd842  : out_data_ref <= 14'h07bf; // 'd1983
      11'd843  : out_data_ref <= 14'h09a2; // 'd2466
      11'd844  : out_data_ref <= 14'h0159; // 'd345
      11'd845  : out_data_ref <= 14'h037e; // 'd894
      11'd846  : out_data_ref <= 14'h0569; // 'd1385
      11'd847  : out_data_ref <= 14'h0884; // 'd2180
      11'd848  : out_data_ref <= 14'h0876; // 'd2166
      11'd849  : out_data_ref <= 14'h0867; // 'd2151
      11'd850  : out_data_ref <= 14'h09eb; // 'd2539
      11'd851  : out_data_ref <= 14'h08a6; // 'd2214
      11'd852  : out_data_ref <= 14'h050e; // 'd1294
      11'd853  : out_data_ref <= 14'h09fc; // 'd2556
      11'd854  : out_data_ref <= 14'h0060; // 'd96
      11'd855  : out_data_ref <= 14'h05ea; // 'd1514
      11'd856  : out_data_ref <= 14'h03d6; // 'd982
      11'd857  : out_data_ref <= 14'h088f; // 'd2191
      11'd858  : out_data_ref <= 14'h03c6; // 'd966
      11'd859  : out_data_ref <= 14'h02e3; // 'd739
      11'd860  : out_data_ref <= 14'h010c; // 'd268
      11'd861  : out_data_ref <= 14'h02ed; // 'd749
      11'd862  : out_data_ref <= 14'h0977; // 'd2423
      11'd863  : out_data_ref <= 14'h09ba; // 'd2490
      11'd864  : out_data_ref <= 14'h0138; // 'd312
      11'd865  : out_data_ref <= 14'h04a5; // 'd1189
      11'd866  : out_data_ref <= 14'h0309; // 'd777
      11'd867  : out_data_ref <= 14'h04b7; // 'd1207
      11'd868  : out_data_ref <= 14'h0898; // 'd2200
      11'd869  : out_data_ref <= 14'h0185; // 'd389
      11'd870  : out_data_ref <= 14'h08d7; // 'd2263
      11'd871  : out_data_ref <= 14'h0446; // 'd1094
      11'd872  : out_data_ref <= 14'h0006; // 'd6
      11'd873  : out_data_ref <= 14'h0679; // 'd1657
      11'd874  : out_data_ref <= 14'h04f2; // 'd1266
      11'd875  : out_data_ref <= 14'h0222; // 'd546
      11'd876  : out_data_ref <= 14'h0144; // 'd324
      11'd877  : out_data_ref <= 14'h02bf; // 'd703
      11'd878  : out_data_ref <= 14'h06e1; // 'd1761
      11'd879  : out_data_ref <= 14'h00c4; // 'd196
      11'd880  : out_data_ref <= 14'h08e4; // 'd2276
      11'd881  : out_data_ref <= 14'h002c; // 'd44
      11'd882  : out_data_ref <= 14'h084f; // 'd2127
      11'd883  : out_data_ref <= 14'h0380; // 'd896
      11'd884  : out_data_ref <= 14'h0494; // 'd1172
      11'd885  : out_data_ref <= 14'h00b5; // 'd181
      11'd886  : out_data_ref <= 14'h0558; // 'd1368
      11'd887  : out_data_ref <= 14'h08e1; // 'd2273
      11'd888  : out_data_ref <= 14'h013e; // 'd318
      11'd889  : out_data_ref <= 14'h05f7; // 'd1527
      11'd890  : out_data_ref <= 14'h03f9; // 'd1017
      11'd891  : out_data_ref <= 14'h00e8; // 'd232
      11'd892  : out_data_ref <= 14'h052f; // 'd1327
      11'd893  : out_data_ref <= 14'h038d; // 'd909
      11'd894  : out_data_ref <= 14'h09ce; // 'd2510
      11'd895  : out_data_ref <= 14'h028e; // 'd654
      11'd896  : out_data_ref <= 14'h0399; // 'd921
      11'd897  : out_data_ref <= 14'h06b1; // 'd1713
      11'd898  : out_data_ref <= 14'h06aa; // 'd1706
      11'd899  : out_data_ref <= 14'h07e3; // 'd2019
      11'd900  : out_data_ref <= 14'h0870; // 'd2160
      11'd901  : out_data_ref <= 14'h00d2; // 'd210
      11'd902  : out_data_ref <= 14'h078d; // 'd1933
      11'd903  : out_data_ref <= 14'h0168; // 'd360
      11'd904  : out_data_ref <= 14'h0229; // 'd553
      11'd905  : out_data_ref <= 14'h014d; // 'd333
      11'd906  : out_data_ref <= 14'h03ec; // 'd1004
      11'd907  : out_data_ref <= 14'h00b7; // 'd183
      11'd908  : out_data_ref <= 14'h0783; // 'd1923
      11'd909  : out_data_ref <= 14'h0745; // 'd1861
      11'd910  : out_data_ref <= 14'h07c8; // 'd1992
      11'd911  : out_data_ref <= 14'h034d; // 'd845
      11'd912  : out_data_ref <= 14'h06fc; // 'd1788
      11'd913  : out_data_ref <= 14'h0470; // 'd1136
      11'd914  : out_data_ref <= 14'h01c7; // 'd455
      11'd915  : out_data_ref <= 14'h0a1b; // 'd2587
      11'd916  : out_data_ref <= 14'h0744; // 'd1860
      11'd917  : out_data_ref <= 14'h06f0; // 'd1776
      11'd918  : out_data_ref <= 14'h033d; // 'd829
      11'd919  : out_data_ref <= 14'h0122; // 'd290
      11'd920  : out_data_ref <= 14'h035c; // 'd860
      11'd921  : out_data_ref <= 14'h0a22; // 'd2594
      11'd922  : out_data_ref <= 14'h0230; // 'd560
      11'd923  : out_data_ref <= 14'h08d5; // 'd2261
      11'd924  : out_data_ref <= 14'h0701; // 'd1793
      11'd925  : out_data_ref <= 14'h0033; // 'd51
      11'd926  : out_data_ref <= 14'h07f9; // 'd2041
      11'd927  : out_data_ref <= 14'h09ff; // 'd2559
      11'd928  : out_data_ref <= 14'h0902; // 'd2306
      11'd929  : out_data_ref <= 14'h033a; // 'd826
      11'd930  : out_data_ref <= 14'h0985; // 'd2437
      11'd931  : out_data_ref <= 14'h0407; // 'd1031
      11'd932  : out_data_ref <= 14'h0736; // 'd1846
      11'd933  : out_data_ref <= 14'h0303; // 'd771
      11'd934  : out_data_ref <= 14'h0460; // 'd1120
      11'd935  : out_data_ref <= 14'h02a4; // 'd676
      11'd936  : out_data_ref <= 14'h0151; // 'd337
      11'd937  : out_data_ref <= 14'h001e; // 'd30
      11'd938  : out_data_ref <= 14'h05b2; // 'd1458
      11'd939  : out_data_ref <= 14'h08d5; // 'd2261
      11'd940  : out_data_ref <= 14'h0869; // 'd2153
      11'd941  : out_data_ref <= 14'h09aa; // 'd2474
      11'd942  : out_data_ref <= 14'h0415; // 'd1045
      11'd943  : out_data_ref <= 14'h07e8; // 'd2024
      11'd944  : out_data_ref <= 14'h034f; // 'd847
      11'd945  : out_data_ref <= 14'h0698; // 'd1688
      11'd946  : out_data_ref <= 14'h09d3; // 'd2515
      11'd947  : out_data_ref <= 14'h058a; // 'd1418
      11'd948  : out_data_ref <= 14'h058e; // 'd1422
      11'd949  : out_data_ref <= 14'h0979; // 'd2425
      11'd950  : out_data_ref <= 14'h0246; // 'd582
      11'd951  : out_data_ref <= 14'h000b; // 'd11
      11'd952  : out_data_ref <= 14'h09ad; // 'd2477
      11'd953  : out_data_ref <= 14'h03b4; // 'd948
      11'd954  : out_data_ref <= 14'h07a6; // 'd1958
      11'd955  : out_data_ref <= 14'h0939; // 'd2361
      11'd956  : out_data_ref <= 14'h0366; // 'd870
      11'd957  : out_data_ref <= 14'h039b; // 'd923
      11'd958  : out_data_ref <= 14'h08dc; // 'd2268
      11'd959  : out_data_ref <= 14'h02f7; // 'd759
      11'd960  : out_data_ref <= 14'h06c7; // 'd1735
      11'd961  : out_data_ref <= 14'h0244; // 'd580
      11'd962  : out_data_ref <= 14'h0569; // 'd1385
      11'd963  : out_data_ref <= 14'h03ae; // 'd942
      11'd964  : out_data_ref <= 14'h086e; // 'd2158
      11'd965  : out_data_ref <= 14'h0182; // 'd386
      11'd966  : out_data_ref <= 14'h06df; // 'd1759
      11'd967  : out_data_ref <= 14'h0923; // 'd2339
      11'd968  : out_data_ref <= 14'h06d2; // 'd1746
      11'd969  : out_data_ref <= 14'h09c5; // 'd2501
      11'd970  : out_data_ref <= 14'h05f8; // 'd1528
      11'd971  : out_data_ref <= 14'h04c6; // 'd1222
      11'd972  : out_data_ref <= 14'h0800; // 'd2048
      11'd973  : out_data_ref <= 14'h0206; // 'd518
      11'd974  : out_data_ref <= 14'h07bb; // 'd1979
      11'd975  : out_data_ref <= 14'h0a33; // 'd2611
      11'd976  : out_data_ref <= 14'h0459; // 'd1113
      11'd977  : out_data_ref <= 14'h039b; // 'd923
      11'd978  : out_data_ref <= 14'h0377; // 'd887
      11'd979  : out_data_ref <= 14'h0921; // 'd2337
      11'd980  : out_data_ref <= 14'h09fc; // 'd2556
      11'd981  : out_data_ref <= 14'h070b; // 'd1803
      11'd982  : out_data_ref <= 14'h0117; // 'd279
      11'd983  : out_data_ref <= 14'h0645; // 'd1605
      11'd984  : out_data_ref <= 14'h0322; // 'd802
      11'd985  : out_data_ref <= 14'h0460; // 'd1120
      11'd986  : out_data_ref <= 14'h073a; // 'd1850
      11'd987  : out_data_ref <= 14'h00e3; // 'd227
      11'd988  : out_data_ref <= 14'h02c3; // 'd707
      11'd989  : out_data_ref <= 14'h0386; // 'd902
      11'd990  : out_data_ref <= 14'h07c6; // 'd1990
      11'd991  : out_data_ref <= 14'h09c0; // 'd2496
      11'd992  : out_data_ref <= 14'h08d7; // 'd2263
      11'd993  : out_data_ref <= 14'h02d4; // 'd724
      11'd994  : out_data_ref <= 14'h0097; // 'd151
      11'd995  : out_data_ref <= 14'h0533; // 'd1331
      11'd996  : out_data_ref <= 14'h08d4; // 'd2260
      11'd997  : out_data_ref <= 14'h070b; // 'd1803
      11'd998  : out_data_ref <= 14'h081a; // 'd2074
      11'd999  : out_data_ref <= 14'h0933; // 'd2355
      11'd1000 : out_data_ref <= 14'h07e7; // 'd2023
      11'd1001 : out_data_ref <= 14'h051a; // 'd1306
      11'd1002 : out_data_ref <= 14'h0393; // 'd915
      11'd1003 : out_data_ref <= 14'h0a0e; // 'd2574
      11'd1004 : out_data_ref <= 14'h08f6; // 'd2294
      11'd1005 : out_data_ref <= 14'h07b9; // 'd1977
      11'd1006 : out_data_ref <= 14'h075f; // 'd1887
      11'd1007 : out_data_ref <= 14'h013c; // 'd316
      11'd1008 : out_data_ref <= 14'h031f; // 'd799
      11'd1009 : out_data_ref <= 14'h021a; // 'd538
      11'd1010 : out_data_ref <= 14'h0287; // 'd647
      11'd1011 : out_data_ref <= 14'h0244; // 'd580
      11'd1012 : out_data_ref <= 14'h0003; // 'd3
      11'd1013 : out_data_ref <= 14'h066d; // 'd1645
      11'd1014 : out_data_ref <= 14'h001c; // 'd28
      11'd1015 : out_data_ref <= 14'h0348; // 'd840
      11'd1016 : out_data_ref <= 14'h026b; // 'd619
      11'd1017 : out_data_ref <= 14'h0161; // 'd353
      11'd1018 : out_data_ref <= 14'h0946; // 'd2374
      11'd1019 : out_data_ref <= 14'h0122; // 'd290
      11'd1020 : out_data_ref <= 14'h05bd; // 'd1469
      11'd1021 : out_data_ref <= 14'h0117; // 'd279
      11'd1022 : out_data_ref <= 14'h04a7; // 'd1191
      11'd1023 : out_data_ref <= 14'h0543; // 'd1347
      11'd1024 : out_data_ref <= 14'h01e2; // 'd482
      11'd1025 : out_data_ref <= 14'h09c9; // 'd2505
      11'd1026 : out_data_ref <= 14'h00d9; // 'd217
      11'd1027 : out_data_ref <= 14'h089e; // 'd2206
      11'd1028 : out_data_ref <= 14'h032c; // 'd812
      11'd1029 : out_data_ref <= 14'h0007; // 'd7
      11'd1030 : out_data_ref <= 14'h0466; // 'd1126
      11'd1031 : out_data_ref <= 14'h0280; // 'd640
      11'd1032 : out_data_ref <= 14'h063f; // 'd1599
      11'd1033 : out_data_ref <= 14'h08cf; // 'd2255
      11'd1034 : out_data_ref <= 14'h0690; // 'd1680
      11'd1035 : out_data_ref <= 14'h073e; // 'd1854
      11'd1036 : out_data_ref <= 14'h09d7; // 'd2519
      11'd1037 : out_data_ref <= 14'h062c; // 'd1580
      11'd1038 : out_data_ref <= 14'h0329; // 'd809
      11'd1039 : out_data_ref <= 14'h02b7; // 'd695
      11'd1040 : out_data_ref <= 14'h0191; // 'd401
      11'd1041 : out_data_ref <= 14'h008c; // 'd140
      11'd1042 : out_data_ref <= 14'h00da; // 'd218
      11'd1043 : out_data_ref <= 14'h0519; // 'd1305
      11'd1044 : out_data_ref <= 14'h01a1; // 'd417
      11'd1045 : out_data_ref <= 14'h05c7; // 'd1479
      11'd1046 : out_data_ref <= 14'h010a; // 'd266
      11'd1047 : out_data_ref <= 14'h06ca; // 'd1738
      11'd1048 : out_data_ref <= 14'h09a8; // 'd2472
      11'd1049 : out_data_ref <= 14'h0667; // 'd1639
      11'd1050 : out_data_ref <= 14'h0885; // 'd2181
      11'd1051 : out_data_ref <= 14'h060a; // 'd1546
      11'd1052 : out_data_ref <= 14'h01f7; // 'd503
      11'd1053 : out_data_ref <= 14'h0902; // 'd2306
      11'd1054 : out_data_ref <= 14'h08a0; // 'd2208
      11'd1055 : out_data_ref <= 14'h0358; // 'd856
      11'd1056 : out_data_ref <= 14'h0347; // 'd839
      11'd1057 : out_data_ref <= 14'h0997; // 'd2455
      11'd1058 : out_data_ref <= 14'h075d; // 'd1885
      11'd1059 : out_data_ref <= 14'h00ad; // 'd173
      11'd1060 : out_data_ref <= 14'h02da; // 'd730
      11'd1061 : out_data_ref <= 14'h094d; // 'd2381
      11'd1062 : out_data_ref <= 14'h00bb; // 'd187
      11'd1063 : out_data_ref <= 14'h0734; // 'd1844
      11'd1064 : out_data_ref <= 14'h0434; // 'd1076
      11'd1065 : out_data_ref <= 14'h06c5; // 'd1733
      11'd1066 : out_data_ref <= 14'h0450; // 'd1104
      11'd1067 : out_data_ref <= 14'h0438; // 'd1080
      11'd1068 : out_data_ref <= 14'h07ad; // 'd1965
      11'd1069 : out_data_ref <= 14'h0531; // 'd1329
      11'd1070 : out_data_ref <= 14'h04a7; // 'd1191
      11'd1071 : out_data_ref <= 14'h0328; // 'd808
      11'd1072 : out_data_ref <= 14'h02f3; // 'd755
      11'd1073 : out_data_ref <= 14'h0181; // 'd385
      11'd1074 : out_data_ref <= 14'h0255; // 'd597
      11'd1075 : out_data_ref <= 14'h012e; // 'd302
      11'd1076 : out_data_ref <= 14'h0525; // 'd1317
      11'd1077 : out_data_ref <= 14'h02bf; // 'd703
      11'd1078 : out_data_ref <= 14'h0131; // 'd305
      11'd1079 : out_data_ref <= 14'h0a34; // 'd2612
      11'd1080 : out_data_ref <= 14'h09f4; // 'd2548
      11'd1081 : out_data_ref <= 14'h0444; // 'd1092
      11'd1082 : out_data_ref <= 14'h089d; // 'd2205
      11'd1083 : out_data_ref <= 14'h05a6; // 'd1446
      11'd1084 : out_data_ref <= 14'h06cc; // 'd1740
      11'd1085 : out_data_ref <= 14'h05b3; // 'd1459
      11'd1086 : out_data_ref <= 14'h07c8; // 'd1992
      11'd1087 : out_data_ref <= 14'h0090; // 'd144
      11'd1088 : out_data_ref <= 14'h09a7; // 'd2471
      11'd1089 : out_data_ref <= 14'h0600; // 'd1536
      11'd1090 : out_data_ref <= 14'h068c; // 'd1676
      11'd1091 : out_data_ref <= 14'h0a2e; // 'd2606
      11'd1092 : out_data_ref <= 14'h016f; // 'd367
      11'd1093 : out_data_ref <= 14'h036f; // 'd879
      11'd1094 : out_data_ref <= 14'h0554; // 'd1364
      11'd1095 : out_data_ref <= 14'h03d4; // 'd980
      11'd1096 : out_data_ref <= 14'h049c; // 'd1180
      11'd1097 : out_data_ref <= 14'h082c; // 'd2092
      11'd1098 : out_data_ref <= 14'h0880; // 'd2176
      11'd1099 : out_data_ref <= 14'h006c; // 'd108
      11'd1100 : out_data_ref <= 14'h03c5; // 'd965
      11'd1101 : out_data_ref <= 14'h09e6; // 'd2534
      11'd1102 : out_data_ref <= 14'h015b; // 'd347
      11'd1103 : out_data_ref <= 14'h061e; // 'd1566
      11'd1104 : out_data_ref <= 14'h0374; // 'd884
      11'd1105 : out_data_ref <= 14'h094c; // 'd2380
      11'd1106 : out_data_ref <= 14'h0827; // 'd2087
      11'd1107 : out_data_ref <= 14'h0593; // 'd1427
      11'd1108 : out_data_ref <= 14'h0042; // 'd66
      11'd1109 : out_data_ref <= 14'h044a; // 'd1098
      11'd1110 : out_data_ref <= 14'h004d; // 'd77
      11'd1111 : out_data_ref <= 14'h04a1; // 'd1185
      11'd1112 : out_data_ref <= 14'h055f; // 'd1375
      11'd1113 : out_data_ref <= 14'h03a0; // 'd928
      11'd1114 : out_data_ref <= 14'h05c0; // 'd1472
      11'd1115 : out_data_ref <= 14'h05f7; // 'd1527
      11'd1116 : out_data_ref <= 14'h0502; // 'd1282
      11'd1117 : out_data_ref <= 14'h06fd; // 'd1789
      11'd1118 : out_data_ref <= 14'h0094; // 'd148
      11'd1119 : out_data_ref <= 14'h0083; // 'd131
      11'd1120 : out_data_ref <= 14'h0957; // 'd2391
      11'd1121 : out_data_ref <= 14'h00a4; // 'd164
      11'd1122 : out_data_ref <= 14'h0230; // 'd560
      11'd1123 : out_data_ref <= 14'h0942; // 'd2370
      11'd1124 : out_data_ref <= 14'h06ed; // 'd1773
      11'd1125 : out_data_ref <= 14'h0320; // 'd800
      11'd1126 : out_data_ref <= 14'h0863; // 'd2147
      11'd1127 : out_data_ref <= 14'h04d1; // 'd1233
      11'd1128 : out_data_ref <= 14'h0951; // 'd2385
      11'd1129 : out_data_ref <= 14'h024d; // 'd589
      11'd1130 : out_data_ref <= 14'h07d9; // 'd2009
      11'd1131 : out_data_ref <= 14'h03e9; // 'd1001
      11'd1132 : out_data_ref <= 14'h0958; // 'd2392
      11'd1133 : out_data_ref <= 14'h034c; // 'd844
      11'd1134 : out_data_ref <= 14'h05d1; // 'd1489
      11'd1135 : out_data_ref <= 14'h08b8; // 'd2232
      11'd1136 : out_data_ref <= 14'h06b0; // 'd1712
      11'd1137 : out_data_ref <= 14'h077b; // 'd1915
      11'd1138 : out_data_ref <= 14'h027a; // 'd634
      11'd1139 : out_data_ref <= 14'h0692; // 'd1682
      11'd1140 : out_data_ref <= 14'h06c0; // 'd1728
      11'd1141 : out_data_ref <= 14'h04e1; // 'd1249
      11'd1142 : out_data_ref <= 14'h0438; // 'd1080
      11'd1143 : out_data_ref <= 14'h01a4; // 'd420
      11'd1144 : out_data_ref <= 14'h030c; // 'd780
      11'd1145 : out_data_ref <= 14'h0761; // 'd1889
      11'd1146 : out_data_ref <= 14'h0920; // 'd2336
      11'd1147 : out_data_ref <= 14'h07e8; // 'd2024
      11'd1148 : out_data_ref <= 14'h0183; // 'd387
      11'd1149 : out_data_ref <= 14'h098e; // 'd2446
      11'd1150 : out_data_ref <= 14'h0681; // 'd1665
      11'd1151 : out_data_ref <= 14'h012c; // 'd300
      11'd1152 : out_data_ref <= 14'h08ab; // 'd2219
      11'd1153 : out_data_ref <= 14'h0022; // 'd34
      11'd1154 : out_data_ref <= 14'h0606; // 'd1542
      11'd1155 : out_data_ref <= 14'h0465; // 'd1125
      11'd1156 : out_data_ref <= 14'h025b; // 'd603
      11'd1157 : out_data_ref <= 14'h08e2; // 'd2274
      11'd1158 : out_data_ref <= 14'h0632; // 'd1586
      11'd1159 : out_data_ref <= 14'h06c7; // 'd1735
      11'd1160 : out_data_ref <= 14'h04e2; // 'd1250
      11'd1161 : out_data_ref <= 14'h000e; // 'd14
      11'd1162 : out_data_ref <= 14'h0a28; // 'd2600
      11'd1163 : out_data_ref <= 14'h04e0; // 'd1248
      11'd1164 : out_data_ref <= 14'h08a2; // 'd2210
      11'd1165 : out_data_ref <= 14'h0650; // 'd1616
      11'd1166 : out_data_ref <= 14'h05d4; // 'd1492
      11'd1167 : out_data_ref <= 14'h096d; // 'd2413
      11'd1168 : out_data_ref <= 14'h08b8; // 'd2232
      11'd1169 : out_data_ref <= 14'h0203; // 'd515
      11'd1170 : out_data_ref <= 14'h0009; // 'd9
      11'd1171 : out_data_ref <= 14'h05ff; // 'd1535
      11'd1172 : out_data_ref <= 14'h045b; // 'd1115
      11'd1173 : out_data_ref <= 14'h0973; // 'd2419
      11'd1174 : out_data_ref <= 14'h05e9; // 'd1513
      11'd1175 : out_data_ref <= 14'h0580; // 'd1408
      11'd1176 : out_data_ref <= 14'h0846; // 'd2118
      11'd1177 : out_data_ref <= 14'h0794; // 'd1940
      11'd1178 : out_data_ref <= 14'h0987; // 'd2439
      11'd1179 : out_data_ref <= 14'h00d9; // 'd217
      11'd1180 : out_data_ref <= 14'h04f4; // 'd1268
      11'd1181 : out_data_ref <= 14'h020e; // 'd526
      11'd1182 : out_data_ref <= 14'h03ca; // 'd970
      11'd1183 : out_data_ref <= 14'h05bf; // 'd1471
      11'd1184 : out_data_ref <= 14'h0871; // 'd2161
      11'd1185 : out_data_ref <= 14'h04d5; // 'd1237
      11'd1186 : out_data_ref <= 14'h077b; // 'd1915
      11'd1187 : out_data_ref <= 14'h053e; // 'd1342
      11'd1188 : out_data_ref <= 14'h04ca; // 'd1226
      11'd1189 : out_data_ref <= 14'h01e5; // 'd485
      11'd1190 : out_data_ref <= 14'h01ca; // 'd458
      11'd1191 : out_data_ref <= 14'h0332; // 'd818
      11'd1192 : out_data_ref <= 14'h04ec; // 'd1260
      11'd1193 : out_data_ref <= 14'h0360; // 'd864
      11'd1194 : out_data_ref <= 14'h04c6; // 'd1222
      11'd1195 : out_data_ref <= 14'h08af; // 'd2223
      11'd1196 : out_data_ref <= 14'h06c5; // 'd1733
      11'd1197 : out_data_ref <= 14'h092b; // 'd2347
      11'd1198 : out_data_ref <= 14'h0649; // 'd1609
      11'd1199 : out_data_ref <= 14'h0355; // 'd853
      11'd1200 : out_data_ref <= 14'h0731; // 'd1841
      11'd1201 : out_data_ref <= 14'h0083; // 'd131
      11'd1202 : out_data_ref <= 14'h02f9; // 'd761
      11'd1203 : out_data_ref <= 14'h074a; // 'd1866
      11'd1204 : out_data_ref <= 14'h0280; // 'd640
      11'd1205 : out_data_ref <= 14'h02be; // 'd702
      11'd1206 : out_data_ref <= 14'h007a; // 'd122
      11'd1207 : out_data_ref <= 14'h043c; // 'd1084
      11'd1208 : out_data_ref <= 14'h0516; // 'd1302
      11'd1209 : out_data_ref <= 14'h054d; // 'd1357
      11'd1210 : out_data_ref <= 14'h0092; // 'd146
      11'd1211 : out_data_ref <= 14'h0863; // 'd2147
      11'd1212 : out_data_ref <= 14'h0910; // 'd2320
      11'd1213 : out_data_ref <= 14'h043a; // 'd1082
      11'd1214 : out_data_ref <= 14'h031b; // 'd795
      11'd1215 : out_data_ref <= 14'h05a9; // 'd1449
      11'd1216 : out_data_ref <= 14'h0a34; // 'd2612
      11'd1217 : out_data_ref <= 14'h01cb; // 'd459
      11'd1218 : out_data_ref <= 14'h02f0; // 'd752
      11'd1219 : out_data_ref <= 14'h04c1; // 'd1217
      11'd1220 : out_data_ref <= 14'h025a; // 'd602
      11'd1221 : out_data_ref <= 14'h04e3; // 'd1251
      11'd1222 : out_data_ref <= 14'h08a5; // 'd2213
      11'd1223 : out_data_ref <= 14'h0993; // 'd2451
      11'd1224 : out_data_ref <= 14'h02de; // 'd734
      11'd1225 : out_data_ref <= 14'h03ae; // 'd942
      11'd1226 : out_data_ref <= 14'h071e; // 'd1822
      11'd1227 : out_data_ref <= 14'h09a9; // 'd2473
      11'd1228 : out_data_ref <= 14'h03c9; // 'd969
      11'd1229 : out_data_ref <= 14'h0126; // 'd294
      11'd1230 : out_data_ref <= 14'h0830; // 'd2096
      11'd1231 : out_data_ref <= 14'h0789; // 'd1929
      11'd1232 : out_data_ref <= 14'h0687; // 'd1671
      11'd1233 : out_data_ref <= 14'h099f; // 'd2463
      11'd1234 : out_data_ref <= 14'h055b; // 'd1371
      11'd1235 : out_data_ref <= 14'h06c6; // 'd1734
      11'd1236 : out_data_ref <= 14'h0118; // 'd280
      11'd1237 : out_data_ref <= 14'h028b; // 'd651
      11'd1238 : out_data_ref <= 14'h08bd; // 'd2237
      11'd1239 : out_data_ref <= 14'h0571; // 'd1393
      11'd1240 : out_data_ref <= 14'h040d; // 'd1037
      11'd1241 : out_data_ref <= 14'h096d; // 'd2413
      11'd1242 : out_data_ref <= 14'h0645; // 'd1605
      11'd1243 : out_data_ref <= 14'h08af; // 'd2223
      11'd1244 : out_data_ref <= 14'h03c5; // 'd965
      11'd1245 : out_data_ref <= 14'h0932; // 'd2354
      11'd1246 : out_data_ref <= 14'h0a29; // 'd2601
      11'd1247 : out_data_ref <= 14'h03e8; // 'd1000
      11'd1248 : out_data_ref <= 14'h03d3; // 'd979
      11'd1249 : out_data_ref <= 14'h08e9; // 'd2281
      11'd1250 : out_data_ref <= 14'h03f9; // 'd1017
      11'd1251 : out_data_ref <= 14'h0475; // 'd1141
      11'd1252 : out_data_ref <= 14'h0957; // 'd2391
      11'd1253 : out_data_ref <= 14'h04fb; // 'd1275
      11'd1254 : out_data_ref <= 14'h0821; // 'd2081
      11'd1255 : out_data_ref <= 14'h07f1; // 'd2033
      11'd1256 : out_data_ref <= 14'h0589; // 'd1417
      11'd1257 : out_data_ref <= 14'h0558; // 'd1368
      11'd1258 : out_data_ref <= 14'h087b; // 'd2171
      11'd1259 : out_data_ref <= 14'h03d3; // 'd979
      11'd1260 : out_data_ref <= 14'h0146; // 'd326
      11'd1261 : out_data_ref <= 14'h0520; // 'd1312
      11'd1262 : out_data_ref <= 14'h01a5; // 'd421
      11'd1263 : out_data_ref <= 14'h005a; // 'd90
      11'd1264 : out_data_ref <= 14'h0373; // 'd883
      11'd1265 : out_data_ref <= 14'h04b9; // 'd1209
      11'd1266 : out_data_ref <= 14'h099c; // 'd2460
      11'd1267 : out_data_ref <= 14'h082d; // 'd2093
      11'd1268 : out_data_ref <= 14'h01d7; // 'd471
      11'd1269 : out_data_ref <= 14'h080d; // 'd2061
      11'd1270 : out_data_ref <= 14'h0823; // 'd2083
      11'd1271 : out_data_ref <= 14'h059b; // 'd1435
      11'd1272 : out_data_ref <= 14'h04e3; // 'd1251
      11'd1273 : out_data_ref <= 14'h0389; // 'd905
      11'd1274 : out_data_ref <= 14'h073a; // 'd1850
      11'd1275 : out_data_ref <= 14'h0506; // 'd1286
      11'd1276 : out_data_ref <= 14'h018a; // 'd394
      default: out_data_ref <= 14'h0;
    endcase
  end

endmodule
