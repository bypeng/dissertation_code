module f_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd1679; // 0
        'h001: dout <=  'sd1595; // 1
        'h002: dout <=  'sd1211; // 2
        'h003: dout <= -'sd1124; // 3
        'h004: dout <= -'sd21; // 4
        'h005: dout <= -'sd232; // 5
        'h006: dout <=  'sd696; // 6
        'h007: dout <=  'sd1326; // 7
        'h008: dout <= -'sd1865; // 8
        'h009: dout <= -'sd2165; // 9
        'h00a: dout <=  'sd1541; // 10
        'h00b: dout <= -'sd309; // 11
        'h00c: dout <=  'sd1204; // 12
        'h00d: dout <= -'sd2286; // 13
        'h00e: dout <= -'sd251; // 14
        'h00f: dout <=  'sd1017; // 15
        'h010: dout <= -'sd1245; // 16
        'h011: dout <=  'sd2044; // 17
        'h012: dout <=  'sd1843; // 18
        'h013: dout <= -'sd2155; // 19
        'h014: dout <= -'sd2179; // 20
        'h015: dout <=  'sd190; // 21
        'h016: dout <=  'sd2016; // 22
        'h017: dout <= -'sd545; // 23
        'h018: dout <= -'sd1301; // 24
        'h019: dout <= -'sd358; // 25
        'h01a: dout <= -'sd2162; // 26
        'h01b: dout <= -'sd1278; // 27
        'h01c: dout <= -'sd285; // 28
        'h01d: dout <= -'sd19; // 29
        'h01e: dout <= -'sd1225; // 30
        'h01f: dout <= -'sd1236; // 31
        'h020: dout <= -'sd1291; // 32
        'h021: dout <= -'sd185; // 33
        'h022: dout <= -'sd965; // 34
        'h023: dout <= -'sd2197; // 35
        'h024: dout <=  'sd1550; // 36
        'h025: dout <=  'sd259; // 37
        'h026: dout <=  'sd653; // 38
        'h027: dout <= -'sd1442; // 39
        'h028: dout <=  'sd2261; // 40
        'h029: dout <=  'sd1653; // 41
        'h02a: dout <= -'sd1740; // 42
        'h02b: dout <= -'sd768; // 43
        'h02c: dout <=  'sd1017; // 44
        'h02d: dout <=  'sd970; // 45
        'h02e: dout <=  'sd2004; // 46
        'h02f: dout <= -'sd358; // 47
        'h030: dout <=  'sd1515; // 48
        'h031: dout <=  'sd782; // 49
        'h032: dout <= -'sd903; // 50
        'h033: dout <=  'sd402; // 51
        'h034: dout <=  'sd1756; // 52
        'h035: dout <=  'sd1589; // 53
        'h036: dout <=  'sd24; // 54
        'h037: dout <=  'sd409; // 55
        'h038: dout <= -'sd2137; // 56
        'h039: dout <= -'sd1181; // 57
        'h03a: dout <=  'sd1365; // 58
        'h03b: dout <= -'sd393; // 59
        'h03c: dout <= -'sd1501; // 60
        'h03d: dout <=  'sd224; // 61
        'h03e: dout <=  'sd932; // 62
        'h03f: dout <=  'sd801; // 63
        'h040: dout <= -'sd575; // 64
        'h041: dout <= -'sd280; // 65
        'h042: dout <=  'sd39; // 66
        'h043: dout <=  'sd1278; // 67
        'h044: dout <=  'sd96; // 68
        'h045: dout <= -'sd490; // 69
        'h046: dout <= -'sd47; // 70
        'h047: dout <= -'sd2160; // 71
        'h048: dout <= -'sd2096; // 72
        'h049: dout <=  'sd934; // 73
        'h04a: dout <=  'sd2218; // 74
        'h04b: dout <=  'sd428; // 75
        'h04c: dout <= -'sd488; // 76
        'h04d: dout <= -'sd1513; // 77
        'h04e: dout <=  'sd10; // 78
        'h04f: dout <=  'sd2213; // 79
        'h050: dout <=  'sd1242; // 80
        'h051: dout <=  'sd182; // 81
        'h052: dout <=  'sd1654; // 82
        'h053: dout <= -'sd1230; // 83
        'h054: dout <=  'sd63; // 84
        'h055: dout <=  'sd2077; // 85
        'h056: dout <=  'sd357; // 86
        'h057: dout <= -'sd188; // 87
        'h058: dout <= -'sd1059; // 88
        'h059: dout <=  'sd220; // 89
        'h05a: dout <=  'sd2099; // 90
        'h05b: dout <= -'sd2269; // 91
        'h05c: dout <=  'sd1302; // 92
        'h05d: dout <=  'sd1471; // 93
        'h05e: dout <=  'sd1773; // 94
        'h05f: dout <=  'sd1104; // 95
        'h060: dout <=  'sd1419; // 96
        'h061: dout <=  'sd86; // 97
        'h062: dout <=  'sd282; // 98
        'h063: dout <= -'sd339; // 99
        'h064: dout <= -'sd2038; // 100
        'h065: dout <=  'sd1699; // 101
        'h066: dout <=  'sd321; // 102
        'h067: dout <= -'sd1378; // 103
        'h068: dout <=  'sd22; // 104
        'h069: dout <= -'sd69; // 105
        'h06a: dout <= -'sd657; // 106
        'h06b: dout <= -'sd707; // 107
        'h06c: dout <=  'sd177; // 108
        'h06d: dout <=  'sd567; // 109
        'h06e: dout <=  'sd516; // 110
        'h06f: dout <= -'sd192; // 111
        'h070: dout <= -'sd2167; // 112
        'h071: dout <= -'sd1241; // 113
        'h072: dout <= -'sd1482; // 114
        'h073: dout <=  'sd388; // 115
        'h074: dout <=  'sd1657; // 116
        'h075: dout <=  'sd1370; // 117
        'h076: dout <=  'sd1364; // 118
        'h077: dout <=  'sd1453; // 119
        'h078: dout <= -'sd1123; // 120
        'h079: dout <=  'sd1569; // 121
        'h07a: dout <=  'sd795; // 122
        'h07b: dout <= -'sd1913; // 123
        'h07c: dout <= -'sd2219; // 124
        'h07d: dout <= -'sd2229; // 125
        'h07e: dout <=  'sd1173; // 126
        'h07f: dout <= -'sd1150; // 127
        'h080: dout <= -'sd1793; // 128
        'h081: dout <=  'sd573; // 129
        'h082: dout <= -'sd714; // 130
        'h083: dout <= -'sd1976; // 131
        'h084: dout <= -'sd1563; // 132
        'h085: dout <=  'sd126; // 133
        'h086: dout <= -'sd1524; // 134
        'h087: dout <= -'sd1043; // 135
        'h088: dout <=  'sd971; // 136
        'h089: dout <= -'sd208; // 137
        'h08a: dout <= -'sd817; // 138
        'h08b: dout <= -'sd120; // 139
        'h08c: dout <= -'sd2187; // 140
        'h08d: dout <= -'sd521; // 141
        'h08e: dout <= -'sd363; // 142
        'h08f: dout <= -'sd1432; // 143
        'h090: dout <= -'sd1796; // 144
        'h091: dout <=  'sd1836; // 145
        'h092: dout <=  'sd46; // 146
        'h093: dout <= -'sd1336; // 147
        'h094: dout <=  'sd485; // 148
        'h095: dout <=  'sd1456; // 149
        'h096: dout <= -'sd2200; // 150
        'h097: dout <= -'sd2213; // 151
        'h098: dout <= -'sd1623; // 152
        'h099: dout <=  'sd1005; // 153
        'h09a: dout <= -'sd1560; // 154
        'h09b: dout <=  'sd939; // 155
        'h09c: dout <=  'sd818; // 156
        'h09d: dout <=  'sd205; // 157
        'h09e: dout <= -'sd1283; // 158
        'h09f: dout <=  'sd2183; // 159
        'h0a0: dout <=  'sd1367; // 160
        'h0a1: dout <=  'sd76; // 161
        'h0a2: dout <= -'sd1271; // 162
        'h0a3: dout <=  'sd682; // 163
        'h0a4: dout <= -'sd483; // 164
        'h0a5: dout <=  'sd348; // 165
        'h0a6: dout <= -'sd821; // 166
        'h0a7: dout <=  'sd601; // 167
        'h0a8: dout <= -'sd2026; // 168
        'h0a9: dout <= -'sd925; // 169
        'h0aa: dout <=  'sd2148; // 170
        'h0ab: dout <=  'sd1724; // 171
        'h0ac: dout <= -'sd889; // 172
        'h0ad: dout <=  'sd1646; // 173
        'h0ae: dout <= -'sd871; // 174
        'h0af: dout <=  'sd2017; // 175
        'h0b0: dout <=  'sd1119; // 176
        'h0b1: dout <= -'sd385; // 177
        'h0b2: dout <= -'sd1137; // 178
        'h0b3: dout <= -'sd2257; // 179
        'h0b4: dout <=  'sd1739; // 180
        'h0b5: dout <= -'sd2121; // 181
        'h0b6: dout <=  'sd1466; // 182
        'h0b7: dout <=  'sd2122; // 183
        'h0b8: dout <=  'sd323; // 184
        'h0b9: dout <= -'sd1508; // 185
        'h0ba: dout <=  'sd1688; // 186
        'h0bb: dout <=  'sd2175; // 187
        'h0bc: dout <=  'sd937; // 188
        'h0bd: dout <=  'sd41; // 189
        'h0be: dout <= -'sd560; // 190
        'h0bf: dout <= -'sd703; // 191
        'h0c0: dout <= -'sd1351; // 192
        'h0c1: dout <=  'sd800; // 193
        'h0c2: dout <= -'sd308; // 194
        'h0c3: dout <= -'sd1404; // 195
        'h0c4: dout <= -'sd1816; // 196
        'h0c5: dout <=  'sd762; // 197
        'h0c6: dout <= -'sd936; // 198
        'h0c7: dout <= -'sd1; // 199
        'h0c8: dout <= -'sd802; // 200
        'h0c9: dout <=  'sd1706; // 201
        'h0ca: dout <=  'sd1835; // 202
        'h0cb: dout <= -'sd2212; // 203
        'h0cc: dout <= -'sd1373; // 204
        'h0cd: dout <= -'sd791; // 205
        'h0ce: dout <=  'sd2236; // 206
        'h0cf: dout <=  'sd1298; // 207
        'h0d0: dout <= -'sd739; // 208
        'h0d1: dout <= -'sd1317; // 209
        'h0d2: dout <=  'sd801; // 210
        'h0d3: dout <=  'sd1550; // 211
        'h0d4: dout <=  'sd1984; // 212
        'h0d5: dout <= -'sd717; // 213
        'h0d6: dout <=  'sd1756; // 214
        'h0d7: dout <=  'sd859; // 215
        'h0d8: dout <= -'sd71; // 216
        'h0d9: dout <=  'sd2229; // 217
        'h0da: dout <= -'sd1218; // 218
        'h0db: dout <=  'sd1035; // 219
        'h0dc: dout <= -'sd1907; // 220
        'h0dd: dout <= -'sd1516; // 221
        'h0de: dout <=  'sd1887; // 222
        'h0df: dout <= -'sd1318; // 223
        'h0e0: dout <=  'sd1190; // 224
        'h0e1: dout <=  'sd460; // 225
        'h0e2: dout <=  'sd1566; // 226
        'h0e3: dout <= -'sd606; // 227
        'h0e4: dout <= -'sd733; // 228
        'h0e5: dout <= -'sd959; // 229
        'h0e6: dout <=  'sd1687; // 230
        'h0e7: dout <=  'sd477; // 231
        'h0e8: dout <=  'sd2086; // 232
        'h0e9: dout <=  'sd1778; // 233
        'h0ea: dout <= -'sd1674; // 234
        'h0eb: dout <=  'sd235; // 235
        'h0ec: dout <= -'sd1817; // 236
        'h0ed: dout <= -'sd2116; // 237
        'h0ee: dout <= -'sd1959; // 238
        'h0ef: dout <=  'sd1681; // 239
        'h0f0: dout <=  'sd1323; // 240
        'h0f1: dout <=  'sd1508; // 241
        'h0f2: dout <= -'sd730; // 242
        'h0f3: dout <=  'sd529; // 243
        'h0f4: dout <=  'sd1294; // 244
        'h0f5: dout <= -'sd560; // 245
        'h0f6: dout <=  'sd325; // 246
        'h0f7: dout <= -'sd1268; // 247
        'h0f8: dout <= -'sd1920; // 248
        'h0f9: dout <= -'sd1071; // 249
        'h0fa: dout <=  'sd1794; // 250
        'h0fb: dout <=  'sd296; // 251
        'h0fc: dout <=  'sd1951; // 252
        'h0fd: dout <= -'sd194; // 253
        'h0fe: dout <= -'sd1023; // 254
        'h0ff: dout <=  'sd1318; // 255
        'h100: dout <=  'sd1505; // 256
        'h101: dout <= -'sd2239; // 257
        'h102: dout <=  'sd782; // 258
        'h103: dout <= -'sd1875; // 259
        'h104: dout <= -'sd1767; // 260
        'h105: dout <=  'sd1768; // 261
        'h106: dout <= -'sd2112; // 262
        'h107: dout <= -'sd1195; // 263
        'h108: dout <=  'sd2241; // 264
        'h109: dout <= -'sd363; // 265
        'h10a: dout <= -'sd1765; // 266
        'h10b: dout <= -'sd1527; // 267
        'h10c: dout <= -'sd1187; // 268
        'h10d: dout <=  'sd1120; // 269
        'h10e: dout <= -'sd1823; // 270
        'h10f: dout <=  'sd1886; // 271
        'h110: dout <= -'sd559; // 272
        'h111: dout <=  'sd2159; // 273
        'h112: dout <=  'sd1879; // 274
        'h113: dout <= -'sd946; // 275
        'h114: dout <= -'sd1132; // 276
        'h115: dout <= -'sd106; // 277
        'h116: dout <= -'sd1836; // 278
        'h117: dout <=  'sd698; // 279
        'h118: dout <= -'sd2114; // 280
        'h119: dout <= -'sd2247; // 281
        'h11a: dout <=  'sd2216; // 282
        'h11b: dout <= -'sd939; // 283
        'h11c: dout <=  'sd443; // 284
        'h11d: dout <= -'sd230; // 285
        'h11e: dout <= -'sd857; // 286
        'h11f: dout <= -'sd2006; // 287
        'h120: dout <=  'sd1898; // 288
        'h121: dout <=  'sd2157; // 289
        'h122: dout <=  'sd2157; // 290
        'h123: dout <= -'sd1784; // 291
        'h124: dout <= -'sd1308; // 292
        'h125: dout <=  'sd541; // 293
        'h126: dout <=  'sd2203; // 294
        'h127: dout <=  'sd197; // 295
        'h128: dout <=  'sd864; // 296
        'h129: dout <=  'sd743; // 297
        'h12a: dout <= -'sd1106; // 298
        'h12b: dout <=  'sd191; // 299
        'h12c: dout <= -'sd885; // 300
        'h12d: dout <= -'sd1164; // 301
        'h12e: dout <= -'sd1922; // 302
        'h12f: dout <= -'sd1006; // 303
        'h130: dout <=  'sd2219; // 304
        'h131: dout <= -'sd239; // 305
        'h132: dout <=  'sd698; // 306
        'h133: dout <=  'sd659; // 307
        'h134: dout <=  'sd2023; // 308
        'h135: dout <= -'sd503; // 309
        'h136: dout <= -'sd887; // 310
        'h137: dout <= -'sd793; // 311
        'h138: dout <= -'sd841; // 312
        'h139: dout <=  'sd1594; // 313
        'h13a: dout <=  'sd1807; // 314
        'h13b: dout <= -'sd905; // 315
        'h13c: dout <= -'sd761; // 316
        'h13d: dout <=  'sd203; // 317
        'h13e: dout <=  'sd363; // 318
        'h13f: dout <=  'sd441; // 319
        'h140: dout <= -'sd1170; // 320
        'h141: dout <= -'sd2202; // 321
        'h142: dout <= -'sd1176; // 322
        'h143: dout <= -'sd1963; // 323
        'h144: dout <=  'sd235; // 324
        'h145: dout <= -'sd1970; // 325
        'h146: dout <= -'sd1951; // 326
        'h147: dout <=  'sd622; // 327
        'h148: dout <= -'sd960; // 328
        'h149: dout <=  'sd1341; // 329
        'h14a: dout <= -'sd31; // 330
        'h14b: dout <=  'sd1665; // 331
        'h14c: dout <= -'sd1588; // 332
        'h14d: dout <=  'sd7; // 333
        'h14e: dout <=  'sd1354; // 334
        'h14f: dout <= -'sd1942; // 335
        'h150: dout <=  'sd2062; // 336
        'h151: dout <= -'sd1500; // 337
        'h152: dout <=  'sd1268; // 338
        'h153: dout <=  'sd2226; // 339
        'h154: dout <=  'sd1476; // 340
        'h155: dout <= -'sd827; // 341
        'h156: dout <= -'sd1805; // 342
        'h157: dout <=  'sd66; // 343
        'h158: dout <=  'sd1925; // 344
        'h159: dout <= -'sd948; // 345
        'h15a: dout <=  'sd1808; // 346
        'h15b: dout <= -'sd1645; // 347
        'h15c: dout <=  'sd1885; // 348
        'h15d: dout <= -'sd2150; // 349
        'h15e: dout <= -'sd844; // 350
        'h15f: dout <=  'sd1851; // 351
        'h160: dout <=  'sd1395; // 352
        'h161: dout <=  'sd1869; // 353
        'h162: dout <=  'sd1564; // 354
        'h163: dout <=  'sd1130; // 355
        'h164: dout <=  'sd870; // 356
        'h165: dout <= -'sd1478; // 357
        'h166: dout <= -'sd309; // 358
        'h167: dout <= -'sd1571; // 359
        'h168: dout <=  'sd986; // 360
        'h169: dout <=  'sd770; // 361
        'h16a: dout <= -'sd1136; // 362
        'h16b: dout <= -'sd2000; // 363
        'h16c: dout <=  'sd2127; // 364
        'h16d: dout <=  'sd1415; // 365
        'h16e: dout <=  'sd226; // 366
        'h16f: dout <=  'sd190; // 367
        'h170: dout <=  'sd1613; // 368
        'h171: dout <= -'sd214; // 369
        'h172: dout <= -'sd479; // 370
        'h173: dout <= -'sd741; // 371
        'h174: dout <= -'sd1111; // 372
        'h175: dout <= -'sd2183; // 373
        'h176: dout <=  'sd672; // 374
        'h177: dout <= -'sd383; // 375
        'h178: dout <=  'sd324; // 376
        'h179: dout <= -'sd2009; // 377
        'h17a: dout <= -'sd666; // 378
        'h17b: dout <= -'sd1661; // 379
        'h17c: dout <= -'sd1721; // 380
        'h17d: dout <= -'sd1106; // 381
        'h17e: dout <=  'sd1510; // 382
        'h17f: dout <= -'sd469; // 383
        'h180: dout <= -'sd454; // 384
        'h181: dout <=  'sd516; // 385
        'h182: dout <= -'sd1223; // 386
        'h183: dout <= -'sd2261; // 387
        'h184: dout <=  'sd132; // 388
        'h185: dout <=  'sd4; // 389
        'h186: dout <=  'sd683; // 390
        'h187: dout <= -'sd283; // 391
        'h188: dout <=  'sd856; // 392
        'h189: dout <=  'sd1062; // 393
        'h18a: dout <= -'sd1201; // 394
        'h18b: dout <= -'sd23; // 395
        'h18c: dout <= -'sd97; // 396
        'h18d: dout <= -'sd1262; // 397
        'h18e: dout <= -'sd403; // 398
        'h18f: dout <=  'sd277; // 399
        'h190: dout <=  'sd1868; // 400
        'h191: dout <=  'sd1918; // 401
        'h192: dout <= -'sd1032; // 402
        'h193: dout <=  'sd672; // 403
        'h194: dout <= -'sd2074; // 404
        'h195: dout <= -'sd1967; // 405
        'h196: dout <=  'sd54; // 406
        'h197: dout <=  'sd1733; // 407
        'h198: dout <= -'sd1563; // 408
        'h199: dout <=  'sd1221; // 409
        'h19a: dout <=  'sd1758; // 410
        'h19b: dout <= -'sd864; // 411
        'h19c: dout <=  'sd884; // 412
        'h19d: dout <=  'sd1602; // 413
        'h19e: dout <= -'sd589; // 414
        'h19f: dout <=  'sd924; // 415
        'h1a0: dout <=  'sd1085; // 416
        'h1a1: dout <=  'sd434; // 417
        'h1a2: dout <=  'sd1636; // 418
        'h1a3: dout <=  'sd1821; // 419
        'h1a4: dout <=  'sd2112; // 420
        'h1a5: dout <=  'sd327; // 421
        'h1a6: dout <= -'sd1486; // 422
        'h1a7: dout <= -'sd1145; // 423
        'h1a8: dout <= -'sd1296; // 424
        'h1a9: dout <=  'sd319; // 425
        'h1aa: dout <=  'sd1183; // 426
        'h1ab: dout <= -'sd2056; // 427
        'h1ac: dout <=  'sd834; // 428
        'h1ad: dout <=  'sd997; // 429
        'h1ae: dout <= -'sd698; // 430
        'h1af: dout <=  'sd69; // 431
        'h1b0: dout <= -'sd1539; // 432
        'h1b1: dout <=  'sd1055; // 433
        'h1b2: dout <= -'sd2109; // 434
        'h1b3: dout <=  'sd2209; // 435
        'h1b4: dout <=  'sd1414; // 436
        'h1b5: dout <=  'sd590; // 437
        'h1b6: dout <= -'sd1067; // 438
        'h1b7: dout <=  'sd1895; // 439
        'h1b8: dout <=  'sd2109; // 440
        'h1b9: dout <= -'sd1657; // 441
        'h1ba: dout <=  'sd1266; // 442
        'h1bb: dout <=  'sd1570; // 443
        'h1bc: dout <=  'sd733; // 444
        'h1bd: dout <=  'sd920; // 445
        'h1be: dout <= -'sd252; // 446
        'h1bf: dout <=  'sd1948; // 447
        'h1c0: dout <=  'sd2163; // 448
        'h1c1: dout <= -'sd540; // 449
        'h1c2: dout <=  'sd1390; // 450
        'h1c3: dout <= -'sd308; // 451
        'h1c4: dout <= -'sd1539; // 452
        'h1c5: dout <= -'sd801; // 453
        'h1c6: dout <= -'sd1716; // 454
        'h1c7: dout <=  'sd1877; // 455
        'h1c8: dout <=  'sd2109; // 456
        'h1c9: dout <= -'sd1748; // 457
        'h1ca: dout <=  'sd462; // 458
        'h1cb: dout <= -'sd421; // 459
        'h1cc: dout <= -'sd1753; // 460
        'h1cd: dout <= -'sd939; // 461
        'h1ce: dout <= -'sd1156; // 462
        'h1cf: dout <=  'sd1146; // 463
        'h1d0: dout <= -'sd2277; // 464
        'h1d1: dout <= -'sd1424; // 465
        'h1d2: dout <= -'sd281; // 466
        'h1d3: dout <= -'sd2199; // 467
        'h1d4: dout <=  'sd585; // 468
        'h1d5: dout <=  'sd485; // 469
        'h1d6: dout <=  'sd1540; // 470
        'h1d7: dout <= -'sd1347; // 471
        'h1d8: dout <= -'sd988; // 472
        'h1d9: dout <=  'sd194; // 473
        'h1da: dout <= -'sd1041; // 474
        'h1db: dout <=  'sd394; // 475
        'h1dc: dout <= -'sd1144; // 476
        'h1dd: dout <=  'sd843; // 477
        'h1de: dout <=  'sd1336; // 478
        'h1df: dout <=  'sd1417; // 479
        'h1e0: dout <=  'sd2174; // 480
        'h1e1: dout <=  'sd208; // 481
        'h1e2: dout <= -'sd42; // 482
        'h1e3: dout <=  'sd1633; // 483
        'h1e4: dout <=  'sd1235; // 484
        'h1e5: dout <=  'sd324; // 485
        'h1e6: dout <= -'sd536; // 486
        'h1e7: dout <= -'sd991; // 487
        'h1e8: dout <= -'sd1799; // 488
        'h1e9: dout <=  'sd1412; // 489
        'h1ea: dout <= -'sd1753; // 490
        'h1eb: dout <=  'sd1135; // 491
        'h1ec: dout <=  'sd208; // 492
        'h1ed: dout <=  'sd2135; // 493
        'h1ee: dout <=  'sd1199; // 494
        'h1ef: dout <=  'sd2174; // 495
        'h1f0: dout <= -'sd1668; // 496
        'h1f1: dout <=  'sd2; // 497
        'h1f2: dout <=  'sd333; // 498
        'h1f3: dout <= -'sd867; // 499
        'h1f4: dout <=  'sd14; // 500
        'h1f5: dout <= -'sd657; // 501
        'h1f6: dout <=  'sd130; // 502
        'h1f7: dout <= -'sd2292; // 503
        'h1f8: dout <= -'sd265; // 504
        'h1f9: dout <= -'sd232; // 505
        'h1fa: dout <= -'sd896; // 506
        'h1fb: dout <= -'sd462; // 507
        'h1fc: dout <=  'sd1300; // 508
        'h1fd: dout <=  'sd842; // 509
        'h1fe: dout <= -'sd35; // 510
        'h1ff: dout <=  'sd678; // 511
        'h200: dout <= -'sd562; // 512
        'h201: dout <= -'sd1359; // 513
        'h202: dout <= -'sd2278; // 514
        'h203: dout <= -'sd1021; // 515
        'h204: dout <=  'sd451; // 516
        'h205: dout <=  'sd1752; // 517
        'h206: dout <=  'sd1512; // 518
        'h207: dout <=  'sd50; // 519
        'h208: dout <=  'sd2236; // 520
        'h209: dout <= -'sd176; // 521
        'h20a: dout <=  'sd1536; // 522
        'h20b: dout <= -'sd418; // 523
        'h20c: dout <=  'sd1123; // 524
        'h20d: dout <=  'sd2239; // 525
        'h20e: dout <= -'sd894; // 526
        'h20f: dout <= -'sd1514; // 527
        'h210: dout <=  'sd551; // 528
        'h211: dout <=  'sd142; // 529
        'h212: dout <= -'sd645; // 530
        'h213: dout <= -'sd2279; // 531
        'h214: dout <= -'sd509; // 532
        'h215: dout <= -'sd340; // 533
        'h216: dout <= -'sd435; // 534
        'h217: dout <=  'sd1658; // 535
        'h218: dout <=  'sd388; // 536
        'h219: dout <=  'sd1074; // 537
        'h21a: dout <=  'sd1827; // 538
        'h21b: dout <=  'sd1142; // 539
        'h21c: dout <= -'sd34; // 540
        'h21d: dout <=  'sd1128; // 541
        'h21e: dout <=  'sd644; // 542
        'h21f: dout <=  'sd683; // 543
        'h220: dout <=  'sd595; // 544
        'h221: dout <= -'sd427; // 545
        'h222: dout <=  'sd593; // 546
        'h223: dout <=  'sd614; // 547
        'h224: dout <=  'sd2007; // 548
        'h225: dout <=  'sd1297; // 549
        'h226: dout <=  'sd1590; // 550
        'h227: dout <=  'sd1228; // 551
        'h228: dout <=  'sd1448; // 552
        'h229: dout <=  'sd484; // 553
        'h22a: dout <= -'sd691; // 554
        'h22b: dout <= -'sd1081; // 555
        'h22c: dout <=  'sd955; // 556
        'h22d: dout <=  'sd1717; // 557
        'h22e: dout <=  'sd203; // 558
        'h22f: dout <= -'sd1597; // 559
        'h230: dout <=  'sd1529; // 560
        'h231: dout <= -'sd71; // 561
        'h232: dout <= -'sd151; // 562
        'h233: dout <= -'sd2087; // 563
        'h234: dout <=  'sd47; // 564
        'h235: dout <=  'sd1124; // 565
        'h236: dout <= -'sd355; // 566
        'h237: dout <= -'sd665; // 567
        'h238: dout <=  'sd720; // 568
        'h239: dout <= -'sd2205; // 569
        'h23a: dout <=  'sd33; // 570
        'h23b: dout <=  'sd2048; // 571
        'h23c: dout <=  'sd874; // 572
        'h23d: dout <= -'sd450; // 573
        'h23e: dout <=  'sd867; // 574
        'h23f: dout <=  'sd482; // 575
        'h240: dout <= -'sd1336; // 576
        'h241: dout <= -'sd1342; // 577
        'h242: dout <=  'sd1772; // 578
        'h243: dout <= -'sd1060; // 579
        'h244: dout <= -'sd1952; // 580
        'h245: dout <=  'sd1518; // 581
        'h246: dout <=  'sd107; // 582
        'h247: dout <= -'sd605; // 583
        'h248: dout <=  'sd53; // 584
        'h249: dout <=  'sd1087; // 585
        'h24a: dout <= -'sd1522; // 586
        'h24b: dout <=  'sd703; // 587
        'h24c: dout <=  'sd980; // 588
        'h24d: dout <=  'sd1446; // 589
        'h24e: dout <= -'sd1057; // 590
        'h24f: dout <=  'sd503; // 591
        'h250: dout <= -'sd1230; // 592
        'h251: dout <=  'sd280; // 593
        'h252: dout <= -'sd1504; // 594
        'h253: dout <=  'sd1330; // 595
        'h254: dout <=  'sd1684; // 596
        'h255: dout <= -'sd782; // 597
        'h256: dout <= -'sd1275; // 598
        'h257: dout <=  'sd2129; // 599
        'h258: dout <=  'sd949; // 600
        'h259: dout <=  'sd1578; // 601
        'h25a: dout <= -'sd2155; // 602
        'h25b: dout <=  'sd1834; // 603
        'h25c: dout <=  'sd562; // 604
        'h25d: dout <= -'sd842; // 605
        'h25e: dout <= -'sd313; // 606
        'h25f: dout <=  'sd1201; // 607
        'h260: dout <=  'sd1310; // 608
        'h261: dout <= -'sd1424; // 609
        'h262: dout <=  'sd578; // 610
        'h263: dout <= -'sd1535; // 611
        'h264: dout <=  'sd2172; // 612
        'h265: dout <= -'sd259; // 613
        'h266: dout <=  'sd1897; // 614
        'h267: dout <=  'sd1048; // 615
        'h268: dout <=  'sd488; // 616
        'h269: dout <= -'sd1093; // 617
        'h26a: dout <=  'sd122; // 618
        'h26b: dout <= -'sd1659; // 619
        'h26c: dout <= -'sd1661; // 620
        'h26d: dout <=  'sd991; // 621
        'h26e: dout <= -'sd638; // 622
        'h26f: dout <=  'sd1154; // 623
        'h270: dout <= -'sd1191; // 624
        'h271: dout <=  'sd1002; // 625
        'h272: dout <=  'sd1003; // 626
        'h273: dout <= -'sd893; // 627
        'h274: dout <= -'sd1807; // 628
        'h275: dout <= -'sd473; // 629
        'h276: dout <= -'sd35; // 630
        'h277: dout <= -'sd1837; // 631
        'h278: dout <= -'sd1438; // 632
        'h279: dout <= -'sd2041; // 633
        'h27a: dout <=  'sd448; // 634
        'h27b: dout <=  'sd1785; // 635
        'h27c: dout <= -'sd1301; // 636
        'h27d: dout <= -'sd2136; // 637
        'h27e: dout <=  'sd936; // 638
        'h27f: dout <=  'sd1446; // 639
        'h280: dout <=  'sd2131; // 640
        'h281: dout <=  'sd520; // 641
        'h282: dout <= -'sd723; // 642
        'h283: dout <=  'sd1551; // 643
        'h284: dout <= -'sd1753; // 644
        'h285: dout <=  'sd884; // 645
        'h286: dout <= -'sd1858; // 646
        'h287: dout <= -'sd460; // 647
        'h288: dout <= -'sd23; // 648
        'h289: dout <= -'sd561; // 649
        'h28a: dout <= -'sd1521; // 650
        'h28b: dout <= -'sd1232; // 651
        'h28c: dout <=  'sd1470; // 652
        'h28d: dout <= -'sd172; // 653
        'h28e: dout <=  'sd367; // 654
        'h28f: dout <= -'sd1323; // 655
        'h290: dout <=  'sd987; // 656
        'h291: dout <= -'sd780; // 657
        'h292: dout <=  'sd430; // 658
        'h293: dout <=  'sd1880; // 659
        'h294: dout <=  'sd2270; // 660
        'h295: dout <= -'sd2083; // 661
        'h296: dout <=  'sd1366; // 662
        'h297: dout <=  'sd1642; // 663
        'h298: dout <= -'sd828; // 664
        'h299: dout <= -'sd536; // 665
        'h29a: dout <=  'sd368; // 666
        'h29b: dout <=  'sd1923; // 667
        'h29c: dout <= -'sd459; // 668
        'h29d: dout <=  'sd1745; // 669
        'h29e: dout <=  'sd1187; // 670
        'h29f: dout <= -'sd1596; // 671
        'h2a0: dout <=  'sd1899; // 672
        'h2a1: dout <= -'sd2226; // 673
        'h2a2: dout <= -'sd1629; // 674
        'h2a3: dout <=  'sd757; // 675
        'h2a4: dout <= -'sd2033; // 676
        'h2a5: dout <= -'sd553; // 677
        'h2a6: dout <= -'sd1699; // 678
        'h2a7: dout <= -'sd170; // 679
        'h2a8: dout <=  'sd1561; // 680
        'h2a9: dout <=  'sd1864; // 681
        'h2aa: dout <= -'sd2133; // 682
        'h2ab: dout <= -'sd2016; // 683
        'h2ac: dout <=  'sd1564; // 684
        'h2ad: dout <= -'sd2099; // 685
        'h2ae: dout <= -'sd1039; // 686
        'h2af: dout <= -'sd1756; // 687
        'h2b0: dout <= -'sd1878; // 688
        'h2b1: dout <= -'sd2169; // 689
        'h2b2: dout <=  'sd631; // 690
        'h2b3: dout <=  'sd1123; // 691
        'h2b4: dout <=  'sd857; // 692
        'h2b5: dout <=  'sd1587; // 693
        'h2b6: dout <=  'sd748; // 694
        'h2b7: dout <= -'sd506; // 695
        'h2b8: dout <=  'sd602; // 696
        'h2b9: dout <=  'sd2156; // 697
        'h2ba: dout <=  'sd650; // 698
        'h2bb: dout <= -'sd1179; // 699
        'h2bc: dout <= -'sd2019; // 700
        'h2bd: dout <=  'sd1998; // 701
        'h2be: dout <=  'sd415; // 702
        'h2bf: dout <= -'sd690; // 703
        'h2c0: dout <=  'sd484; // 704
        'h2c1: dout <=  'sd277; // 705
        'h2c2: dout <=  'sd102; // 706
        'h2c3: dout <= -'sd2016; // 707
        'h2c4: dout <= -'sd674; // 708
        'h2c5: dout <= -'sd401; // 709
        'h2c6: dout <= -'sd1380; // 710
        'h2c7: dout <=  'sd1745; // 711
        'h2c8: dout <= -'sd348; // 712
        'h2c9: dout <=  'sd746; // 713
        'h2ca: dout <=  'sd980; // 714
        'h2cb: dout <=  'sd1117; // 715
        'h2cc: dout <=  'sd1015; // 716
        'h2cd: dout <=  'sd1158; // 717
        'h2ce: dout <= -'sd1140; // 718
        'h2cf: dout <=  'sd2187; // 719
        'h2d0: dout <= -'sd1602; // 720
        'h2d1: dout <=  'sd1922; // 721
        'h2d2: dout <=  'sd1628; // 722
        'h2d3: dout <=  'sd1617; // 723
        'h2d4: dout <= -'sd2053; // 724
        'h2d5: dout <= -'sd1877; // 725
        'h2d6: dout <=  'sd1437; // 726
        'h2d7: dout <= -'sd142; // 727
        'h2d8: dout <= -'sd596; // 728
        'h2d9: dout <=  'sd2225; // 729
        'h2da: dout <= -'sd2111; // 730
        'h2db: dout <=  'sd144; // 731
        'h2dc: dout <= -'sd260; // 732
        'h2dd: dout <= -'sd1707; // 733
        'h2de: dout <= -'sd481; // 734
        'h2df: dout <=  'sd953; // 735
        'h2e0: dout <=  'sd1755; // 736
        'h2e1: dout <= -'sd2182; // 737
        'h2e2: dout <=  'sd113; // 738
        'h2e3: dout <= -'sd1881; // 739
        'h2e4: dout <=  'sd1379; // 740
        'h2e5: dout <= -'sd1902; // 741
        'h2e6: dout <= -'sd2139; // 742
        'h2e7: dout <= -'sd531; // 743
        'h2e8: dout <=  'sd1068; // 744
        'h2e9: dout <= -'sd858; // 745
        'h2ea: dout <= -'sd1699; // 746
        'h2eb: dout <=  'sd1352; // 747
        'h2ec: dout <=  'sd1409; // 748
        'h2ed: dout <=  'sd1634; // 749
        'h2ee: dout <= -'sd901; // 750
        'h2ef: dout <= -'sd345; // 751
        'h2f0: dout <= -'sd1169; // 752
        'h2f1: dout <=  'sd263; // 753
        'h2f2: dout <= -'sd780; // 754
        'h2f3: dout <= -'sd741; // 755
        'h2f4: dout <=  'sd1302; // 756
        'h2f5: dout <=  'sd2095; // 757
        'h2f6: dout <=  'sd386; // 758
        'h2f7: dout <= -'sd1815; // 759
        'h2f8: dout <=  'sd700; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module g_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd236; // 0
        'h001: dout <=  'sd2241; // 1
        'h002: dout <=  'sd1007; // 2
        'h003: dout <=  'sd1537; // 3
        'h004: dout <=  'sd924; // 4
        'h005: dout <=  'sd164; // 5
        'h006: dout <=  'sd1822; // 6
        'h007: dout <=  'sd1522; // 7
        'h008: dout <= -'sd958; // 8
        'h009: dout <= -'sd1575; // 9
        'h00a: dout <= -'sd595; // 10
        'h00b: dout <=  'sd97; // 11
        'h00c: dout <= -'sd1848; // 12
        'h00d: dout <= -'sd710; // 13
        'h00e: dout <=  'sd344; // 14
        'h00f: dout <= -'sd2095; // 15
        'h010: dout <=  'sd1446; // 16
        'h011: dout <=  'sd694; // 17
        'h012: dout <= -'sd856; // 18
        'h013: dout <= -'sd926; // 19
        'h014: dout <= -'sd677; // 20
        'h015: dout <= -'sd802; // 21
        'h016: dout <=  'sd1141; // 22
        'h017: dout <=  'sd5; // 23
        'h018: dout <=  'sd120; // 24
        'h019: dout <= -'sd1613; // 25
        'h01a: dout <=  'sd1903; // 26
        'h01b: dout <= -'sd801; // 27
        'h01c: dout <= -'sd792; // 28
        'h01d: dout <= -'sd1979; // 29
        'h01e: dout <=  'sd2201; // 30
        'h01f: dout <= -'sd93; // 31
        'h020: dout <=  'sd1896; // 32
        'h021: dout <=  'sd1963; // 33
        'h022: dout <=  'sd2157; // 34
        'h023: dout <=  'sd1449; // 35
        'h024: dout <=  'sd1953; // 36
        'h025: dout <=  'sd1939; // 37
        'h026: dout <=  'sd1384; // 38
        'h027: dout <= -'sd1678; // 39
        'h028: dout <=  'sd109; // 40
        'h029: dout <=  'sd347; // 41
        'h02a: dout <=  'sd2261; // 42
        'h02b: dout <=  'sd1304; // 43
        'h02c: dout <=  'sd932; // 44
        'h02d: dout <=  'sd1132; // 45
        'h02e: dout <= -'sd635; // 46
        'h02f: dout <=  'sd2031; // 47
        'h030: dout <=  'sd659; // 48
        'h031: dout <= -'sd447; // 49
        'h032: dout <= -'sd163; // 50
        'h033: dout <=  'sd2203; // 51
        'h034: dout <=  'sd148; // 52
        'h035: dout <= -'sd1525; // 53
        'h036: dout <= -'sd1614; // 54
        'h037: dout <=  'sd860; // 55
        'h038: dout <=  'sd288; // 56
        'h039: dout <=  'sd1868; // 57
        'h03a: dout <= -'sd1448; // 58
        'h03b: dout <= -'sd408; // 59
        'h03c: dout <=  'sd1047; // 60
        'h03d: dout <= -'sd2065; // 61
        'h03e: dout <= -'sd1840; // 62
        'h03f: dout <=  'sd210; // 63
        'h040: dout <= -'sd1076; // 64
        'h041: dout <= -'sd1805; // 65
        'h042: dout <= -'sd1094; // 66
        'h043: dout <=  'sd607; // 67
        'h044: dout <=  'sd121; // 68
        'h045: dout <= -'sd1935; // 69
        'h046: dout <= -'sd1961; // 70
        'h047: dout <=  'sd1610; // 71
        'h048: dout <=  'sd658; // 72
        'h049: dout <= -'sd1500; // 73
        'h04a: dout <=  'sd1661; // 74
        'h04b: dout <= -'sd2195; // 75
        'h04c: dout <= -'sd606; // 76
        'h04d: dout <=  'sd1596; // 77
        'h04e: dout <=  'sd965; // 78
        'h04f: dout <= -'sd993; // 79
        'h050: dout <=  'sd1796; // 80
        'h051: dout <=  'sd450; // 81
        'h052: dout <=  'sd1678; // 82
        'h053: dout <=  'sd1803; // 83
        'h054: dout <= -'sd342; // 84
        'h055: dout <=  'sd806; // 85
        'h056: dout <=  'sd204; // 86
        'h057: dout <=  'sd2042; // 87
        'h058: dout <=  'sd1369; // 88
        'h059: dout <=  'sd1037; // 89
        'h05a: dout <=  'sd1442; // 90
        'h05b: dout <=  'sd2287; // 91
        'h05c: dout <= -'sd1118; // 92
        'h05d: dout <= -'sd1371; // 93
        'h05e: dout <=  'sd1133; // 94
        'h05f: dout <=  'sd1241; // 95
        'h060: dout <=  'sd66; // 96
        'h061: dout <= -'sd59; // 97
        'h062: dout <= -'sd442; // 98
        'h063: dout <=  'sd1757; // 99
        'h064: dout <=  'sd1360; // 100
        'h065: dout <=  'sd388; // 101
        'h066: dout <= -'sd2111; // 102
        'h067: dout <=  'sd1612; // 103
        'h068: dout <= -'sd191; // 104
        'h069: dout <= -'sd1424; // 105
        'h06a: dout <= -'sd921; // 106
        'h06b: dout <=  'sd878; // 107
        'h06c: dout <= -'sd2270; // 108
        'h06d: dout <= -'sd1744; // 109
        'h06e: dout <= -'sd906; // 110
        'h06f: dout <=  'sd1778; // 111
        'h070: dout <=  'sd1133; // 112
        'h071: dout <=  'sd2161; // 113
        'h072: dout <=  'sd198; // 114
        'h073: dout <=  'sd330; // 115
        'h074: dout <=  'sd236; // 116
        'h075: dout <=  'sd118; // 117
        'h076: dout <=  'sd193; // 118
        'h077: dout <=  'sd1463; // 119
        'h078: dout <=  'sd2081; // 120
        'h079: dout <= -'sd421; // 121
        'h07a: dout <=  'sd597; // 122
        'h07b: dout <= -'sd883; // 123
        'h07c: dout <= -'sd909; // 124
        'h07d: dout <=  'sd29; // 125
        'h07e: dout <=  'sd396; // 126
        'h07f: dout <=  'sd230; // 127
        'h080: dout <=  'sd2188; // 128
        'h081: dout <= -'sd1547; // 129
        'h082: dout <=  'sd627; // 130
        'h083: dout <=  'sd2270; // 131
        'h084: dout <=  'sd1084; // 132
        'h085: dout <=  'sd303; // 133
        'h086: dout <= -'sd604; // 134
        'h087: dout <= -'sd449; // 135
        'h088: dout <=  'sd2004; // 136
        'h089: dout <=  'sd1815; // 137
        'h08a: dout <=  'sd779; // 138
        'h08b: dout <=  'sd1831; // 139
        'h08c: dout <=  'sd1952; // 140
        'h08d: dout <=  'sd1590; // 141
        'h08e: dout <= -'sd535; // 142
        'h08f: dout <= -'sd164; // 143
        'h090: dout <=  'sd1359; // 144
        'h091: dout <= -'sd585; // 145
        'h092: dout <=  'sd1145; // 146
        'h093: dout <= -'sd85; // 147
        'h094: dout <= -'sd750; // 148
        'h095: dout <= -'sd201; // 149
        'h096: dout <= -'sd1761; // 150
        'h097: dout <= -'sd668; // 151
        'h098: dout <= -'sd389; // 152
        'h099: dout <= -'sd2212; // 153
        'h09a: dout <= -'sd1506; // 154
        'h09b: dout <= -'sd1101; // 155
        'h09c: dout <=  'sd1643; // 156
        'h09d: dout <=  'sd411; // 157
        'h09e: dout <= -'sd977; // 158
        'h09f: dout <=  'sd2285; // 159
        'h0a0: dout <= -'sd1111; // 160
        'h0a1: dout <=  'sd63; // 161
        'h0a2: dout <=  'sd1100; // 162
        'h0a3: dout <=  'sd878; // 163
        'h0a4: dout <= -'sd305; // 164
        'h0a5: dout <=  'sd1272; // 165
        'h0a6: dout <= -'sd65; // 166
        'h0a7: dout <=  'sd989; // 167
        'h0a8: dout <= -'sd40; // 168
        'h0a9: dout <=  'sd2165; // 169
        'h0aa: dout <=  'sd992; // 170
        'h0ab: dout <= -'sd1876; // 171
        'h0ac: dout <= -'sd1701; // 172
        'h0ad: dout <=  'sd2142; // 173
        'h0ae: dout <= -'sd1243; // 174
        'h0af: dout <= -'sd2176; // 175
        'h0b0: dout <= -'sd1133; // 176
        'h0b1: dout <= -'sd93; // 177
        'h0b2: dout <=  'sd2076; // 178
        'h0b3: dout <= -'sd463; // 179
        'h0b4: dout <=  'sd1026; // 180
        'h0b5: dout <=  'sd1535; // 181
        'h0b6: dout <= -'sd1886; // 182
        'h0b7: dout <=  'sd514; // 183
        'h0b8: dout <=  'sd2276; // 184
        'h0b9: dout <=  'sd228; // 185
        'h0ba: dout <=  'sd158; // 186
        'h0bb: dout <= -'sd704; // 187
        'h0bc: dout <=  'sd2048; // 188
        'h0bd: dout <=  'sd2156; // 189
        'h0be: dout <= -'sd1822; // 190
        'h0bf: dout <=  'sd243; // 191
        'h0c0: dout <= -'sd369; // 192
        'h0c1: dout <=  'sd788; // 193
        'h0c2: dout <= -'sd1751; // 194
        'h0c3: dout <= -'sd1077; // 195
        'h0c4: dout <= -'sd1016; // 196
        'h0c5: dout <= -'sd93; // 197
        'h0c6: dout <=  'sd1346; // 198
        'h0c7: dout <=  'sd1643; // 199
        'h0c8: dout <=  'sd1315; // 200
        'h0c9: dout <=  'sd812; // 201
        'h0ca: dout <= -'sd1895; // 202
        'h0cb: dout <= -'sd506; // 203
        'h0cc: dout <=  'sd775; // 204
        'h0cd: dout <= -'sd945; // 205
        'h0ce: dout <=  'sd36; // 206
        'h0cf: dout <=  'sd1860; // 207
        'h0d0: dout <= -'sd1762; // 208
        'h0d1: dout <=  'sd1625; // 209
        'h0d2: dout <= -'sd1810; // 210
        'h0d3: dout <= -'sd522; // 211
        'h0d4: dout <=  'sd1861; // 212
        'h0d5: dout <= -'sd1372; // 213
        'h0d6: dout <=  'sd95; // 214
        'h0d7: dout <= -'sd383; // 215
        'h0d8: dout <=  'sd1781; // 216
        'h0d9: dout <=  'sd2259; // 217
        'h0da: dout <= -'sd971; // 218
        'h0db: dout <= -'sd35; // 219
        'h0dc: dout <=  'sd1813; // 220
        'h0dd: dout <=  'sd206; // 221
        'h0de: dout <= -'sd1310; // 222
        'h0df: dout <=  'sd1192; // 223
        'h0e0: dout <= -'sd748; // 224
        'h0e1: dout <= -'sd64; // 225
        'h0e2: dout <= -'sd2256; // 226
        'h0e3: dout <=  'sd2245; // 227
        'h0e4: dout <=  'sd722; // 228
        'h0e5: dout <=  'sd1955; // 229
        'h0e6: dout <=  'sd2152; // 230
        'h0e7: dout <= -'sd1067; // 231
        'h0e8: dout <=  'sd186; // 232
        'h0e9: dout <= -'sd274; // 233
        'h0ea: dout <=  'sd1193; // 234
        'h0eb: dout <=  'sd1572; // 235
        'h0ec: dout <= -'sd1246; // 236
        'h0ed: dout <= -'sd1035; // 237
        'h0ee: dout <=  'sd947; // 238
        'h0ef: dout <= -'sd406; // 239
        'h0f0: dout <= -'sd1698; // 240
        'h0f1: dout <= -'sd1399; // 241
        'h0f2: dout <=  'sd279; // 242
        'h0f3: dout <=  'sd452; // 243
        'h0f4: dout <=  'sd2112; // 244
        'h0f5: dout <=  'sd150; // 245
        'h0f6: dout <=  'sd500; // 246
        'h0f7: dout <= -'sd1612; // 247
        'h0f8: dout <= -'sd396; // 248
        'h0f9: dout <= -'sd1011; // 249
        'h0fa: dout <=  'sd897; // 250
        'h0fb: dout <= -'sd1069; // 251
        'h0fc: dout <= -'sd1311; // 252
        'h0fd: dout <= -'sd607; // 253
        'h0fe: dout <= -'sd135; // 254
        'h0ff: dout <= -'sd742; // 255
        'h100: dout <=  'sd485; // 256
        'h101: dout <= -'sd1464; // 257
        'h102: dout <=  'sd1744; // 258
        'h103: dout <=  'sd891; // 259
        'h104: dout <=  'sd160; // 260
        'h105: dout <= -'sd2028; // 261
        'h106: dout <= -'sd799; // 262
        'h107: dout <=  'sd873; // 263
        'h108: dout <=  'sd666; // 264
        'h109: dout <=  'sd1432; // 265
        'h10a: dout <=  'sd1797; // 266
        'h10b: dout <= -'sd848; // 267
        'h10c: dout <= -'sd29; // 268
        'h10d: dout <= -'sd780; // 269
        'h10e: dout <= -'sd1708; // 270
        'h10f: dout <= -'sd1652; // 271
        'h110: dout <= -'sd1118; // 272
        'h111: dout <= -'sd1891; // 273
        'h112: dout <=  'sd178; // 274
        'h113: dout <=  'sd932; // 275
        'h114: dout <=  'sd290; // 276
        'h115: dout <=  'sd848; // 277
        'h116: dout <= -'sd1257; // 278
        'h117: dout <= -'sd1380; // 279
        'h118: dout <=  'sd310; // 280
        'h119: dout <=  'sd1764; // 281
        'h11a: dout <= -'sd357; // 282
        'h11b: dout <= -'sd2276; // 283
        'h11c: dout <= -'sd2203; // 284
        'h11d: dout <= -'sd894; // 285
        'h11e: dout <=  'sd530; // 286
        'h11f: dout <= -'sd1907; // 287
        'h120: dout <= -'sd1265; // 288
        'h121: dout <=  'sd830; // 289
        'h122: dout <=  'sd2227; // 290
        'h123: dout <= -'sd730; // 291
        'h124: dout <=  'sd464; // 292
        'h125: dout <=  'sd85; // 293
        'h126: dout <= -'sd2189; // 294
        'h127: dout <= -'sd781; // 295
        'h128: dout <= -'sd1655; // 296
        'h129: dout <= -'sd1144; // 297
        'h12a: dout <=  'sd1239; // 298
        'h12b: dout <=  'sd832; // 299
        'h12c: dout <= -'sd2107; // 300
        'h12d: dout <= -'sd1940; // 301
        'h12e: dout <=  'sd1033; // 302
        'h12f: dout <= -'sd1822; // 303
        'h130: dout <= -'sd840; // 304
        'h131: dout <= -'sd1059; // 305
        'h132: dout <= -'sd2067; // 306
        'h133: dout <= -'sd2152; // 307
        'h134: dout <= -'sd1657; // 308
        'h135: dout <= -'sd462; // 309
        'h136: dout <=  'sd1991; // 310
        'h137: dout <=  'sd635; // 311
        'h138: dout <= -'sd1184; // 312
        'h139: dout <=  'sd825; // 313
        'h13a: dout <= -'sd1039; // 314
        'h13b: dout <=  'sd70; // 315
        'h13c: dout <= -'sd818; // 316
        'h13d: dout <=  'sd2060; // 317
        'h13e: dout <= -'sd678; // 318
        'h13f: dout <=  'sd1394; // 319
        'h140: dout <=  'sd648; // 320
        'h141: dout <=  'sd1576; // 321
        'h142: dout <=  'sd487; // 322
        'h143: dout <=  'sd1700; // 323
        'h144: dout <= -'sd435; // 324
        'h145: dout <=  'sd822; // 325
        'h146: dout <=  'sd554; // 326
        'h147: dout <=  'sd127; // 327
        'h148: dout <=  'sd296; // 328
        'h149: dout <=  'sd164; // 329
        'h14a: dout <= -'sd488; // 330
        'h14b: dout <=  'sd1829; // 331
        'h14c: dout <=  'sd609; // 332
        'h14d: dout <=  'sd226; // 333
        'h14e: dout <= -'sd2048; // 334
        'h14f: dout <=  'sd39; // 335
        'h150: dout <= -'sd1491; // 336
        'h151: dout <= -'sd1308; // 337
        'h152: dout <= -'sd300; // 338
        'h153: dout <=  'sd211; // 339
        'h154: dout <= -'sd1146; // 340
        'h155: dout <= -'sd1052; // 341
        'h156: dout <=  'sd138; // 342
        'h157: dout <= -'sd123; // 343
        'h158: dout <= -'sd444; // 344
        'h159: dout <= -'sd1819; // 345
        'h15a: dout <= -'sd581; // 346
        'h15b: dout <=  'sd709; // 347
        'h15c: dout <=  'sd203; // 348
        'h15d: dout <=  'sd205; // 349
        'h15e: dout <=  'sd1578; // 350
        'h15f: dout <=  'sd1025; // 351
        'h160: dout <=  'sd847; // 352
        'h161: dout <= -'sd2156; // 353
        'h162: dout <= -'sd881; // 354
        'h163: dout <=  'sd837; // 355
        'h164: dout <= -'sd1580; // 356
        'h165: dout <=  'sd1898; // 357
        'h166: dout <= -'sd1644; // 358
        'h167: dout <=  'sd1741; // 359
        'h168: dout <= -'sd1303; // 360
        'h169: dout <=  'sd1568; // 361
        'h16a: dout <=  'sd1599; // 362
        'h16b: dout <= -'sd755; // 363
        'h16c: dout <=  'sd1784; // 364
        'h16d: dout <= -'sd1562; // 365
        'h16e: dout <=  'sd1603; // 366
        'h16f: dout <= -'sd543; // 367
        'h170: dout <= -'sd277; // 368
        'h171: dout <= -'sd1754; // 369
        'h172: dout <=  'sd464; // 370
        'h173: dout <= -'sd1057; // 371
        'h174: dout <=  'sd766; // 372
        'h175: dout <=  'sd1374; // 373
        'h176: dout <=  'sd476; // 374
        'h177: dout <= -'sd2258; // 375
        'h178: dout <=  'sd2077; // 376
        'h179: dout <=  'sd1927; // 377
        'h17a: dout <=  'sd656; // 378
        'h17b: dout <= -'sd553; // 379
        'h17c: dout <=  'sd284; // 380
        'h17d: dout <=  'sd1757; // 381
        'h17e: dout <= -'sd186; // 382
        'h17f: dout <=  'sd1282; // 383
        'h180: dout <=  'sd452; // 384
        'h181: dout <= -'sd357; // 385
        'h182: dout <=  'sd1990; // 386
        'h183: dout <= -'sd420; // 387
        'h184: dout <=  'sd486; // 388
        'h185: dout <= -'sd2051; // 389
        'h186: dout <= -'sd134; // 390
        'h187: dout <= -'sd2124; // 391
        'h188: dout <=  'sd937; // 392
        'h189: dout <= -'sd2293; // 393
        'h18a: dout <= -'sd2102; // 394
        'h18b: dout <= -'sd1785; // 395
        'h18c: dout <= -'sd1655; // 396
        'h18d: dout <=  'sd37; // 397
        'h18e: dout <= -'sd660; // 398
        'h18f: dout <= -'sd1052; // 399
        'h190: dout <=  'sd2220; // 400
        'h191: dout <=  'sd1878; // 401
        'h192: dout <=  'sd711; // 402
        'h193: dout <=  'sd1387; // 403
        'h194: dout <=  'sd1468; // 404
        'h195: dout <= -'sd1170; // 405
        'h196: dout <=  'sd1415; // 406
        'h197: dout <= -'sd1195; // 407
        'h198: dout <=  'sd286; // 408
        'h199: dout <= -'sd653; // 409
        'h19a: dout <= -'sd1567; // 410
        'h19b: dout <=  'sd1271; // 411
        'h19c: dout <=  'sd1911; // 412
        'h19d: dout <= -'sd855; // 413
        'h19e: dout <=  'sd1743; // 414
        'h19f: dout <= -'sd706; // 415
        'h1a0: dout <=  'sd723; // 416
        'h1a1: dout <=  'sd2276; // 417
        'h1a2: dout <=  'sd1249; // 418
        'h1a3: dout <= -'sd2040; // 419
        'h1a4: dout <= -'sd299; // 420
        'h1a5: dout <= -'sd568; // 421
        'h1a6: dout <= -'sd946; // 422
        'h1a7: dout <=  'sd1451; // 423
        'h1a8: dout <= -'sd271; // 424
        'h1a9: dout <=  'sd915; // 425
        'h1aa: dout <=  'sd619; // 426
        'h1ab: dout <=  'sd87; // 427
        'h1ac: dout <= -'sd2038; // 428
        'h1ad: dout <=  'sd794; // 429
        'h1ae: dout <=  'sd1797; // 430
        'h1af: dout <= -'sd1505; // 431
        'h1b0: dout <=  'sd655; // 432
        'h1b1: dout <= -'sd58; // 433
        'h1b2: dout <= -'sd730; // 434
        'h1b3: dout <=  'sd966; // 435
        'h1b4: dout <=  'sd2182; // 436
        'h1b5: dout <= -'sd2196; // 437
        'h1b6: dout <=  'sd1824; // 438
        'h1b7: dout <= -'sd536; // 439
        'h1b8: dout <=  'sd1533; // 440
        'h1b9: dout <= -'sd1493; // 441
        'h1ba: dout <=  'sd994; // 442
        'h1bb: dout <= -'sd1838; // 443
        'h1bc: dout <= -'sd755; // 444
        'h1bd: dout <=  'sd2157; // 445
        'h1be: dout <=  'sd719; // 446
        'h1bf: dout <=  'sd1306; // 447
        'h1c0: dout <= -'sd178; // 448
        'h1c1: dout <= -'sd132; // 449
        'h1c2: dout <= -'sd34; // 450
        'h1c3: dout <=  'sd1254; // 451
        'h1c4: dout <=  'sd1025; // 452
        'h1c5: dout <= -'sd1406; // 453
        'h1c6: dout <= -'sd273; // 454
        'h1c7: dout <=  'sd193; // 455
        'h1c8: dout <=  'sd328; // 456
        'h1c9: dout <=  'sd1959; // 457
        'h1ca: dout <=  'sd1560; // 458
        'h1cb: dout <= -'sd1607; // 459
        'h1cc: dout <= -'sd569; // 460
        'h1cd: dout <= -'sd1795; // 461
        'h1ce: dout <= -'sd2175; // 462
        'h1cf: dout <= -'sd1953; // 463
        'h1d0: dout <= -'sd1456; // 464
        'h1d1: dout <=  'sd1222; // 465
        'h1d2: dout <=  'sd768; // 466
        'h1d3: dout <=  'sd1368; // 467
        'h1d4: dout <= -'sd971; // 468
        'h1d5: dout <= -'sd1582; // 469
        'h1d6: dout <=  'sd2167; // 470
        'h1d7: dout <=  'sd1497; // 471
        'h1d8: dout <=  'sd2051; // 472
        'h1d9: dout <= -'sd2209; // 473
        'h1da: dout <= -'sd475; // 474
        'h1db: dout <=  'sd614; // 475
        'h1dc: dout <=  'sd1084; // 476
        'h1dd: dout <=  'sd1894; // 477
        'h1de: dout <=  'sd173; // 478
        'h1df: dout <= -'sd501; // 479
        'h1e0: dout <= -'sd2271; // 480
        'h1e1: dout <=  'sd1395; // 481
        'h1e2: dout <=  'sd2214; // 482
        'h1e3: dout <=  'sd1870; // 483
        'h1e4: dout <=  'sd745; // 484
        'h1e5: dout <= -'sd723; // 485
        'h1e6: dout <= -'sd1198; // 486
        'h1e7: dout <=  'sd1263; // 487
        'h1e8: dout <=  'sd1999; // 488
        'h1e9: dout <=  'sd2113; // 489
        'h1ea: dout <= -'sd1489; // 490
        'h1eb: dout <=  'sd392; // 491
        'h1ec: dout <=  'sd60; // 492
        'h1ed: dout <= -'sd333; // 493
        'h1ee: dout <=  'sd1352; // 494
        'h1ef: dout <=  'sd2001; // 495
        'h1f0: dout <=  'sd1031; // 496
        'h1f1: dout <=  'sd920; // 497
        'h1f2: dout <=  'sd875; // 498
        'h1f3: dout <=  'sd705; // 499
        'h1f4: dout <=  'sd169; // 500
        'h1f5: dout <= -'sd1157; // 501
        'h1f6: dout <=  'sd1283; // 502
        'h1f7: dout <= -'sd1749; // 503
        'h1f8: dout <=  'sd661; // 504
        'h1f9: dout <= -'sd519; // 505
        'h1fa: dout <=  'sd275; // 506
        'h1fb: dout <=  'sd649; // 507
        'h1fc: dout <= -'sd97; // 508
        'h1fd: dout <=  'sd2195; // 509
        'h1fe: dout <= -'sd1197; // 510
        'h1ff: dout <= -'sd2240; // 511
        'h200: dout <=  'sd2090; // 512
        'h201: dout <= -'sd863; // 513
        'h202: dout <= -'sd1019; // 514
        'h203: dout <= -'sd388; // 515
        'h204: dout <=  'sd436; // 516
        'h205: dout <=  'sd2232; // 517
        'h206: dout <=  'sd953; // 518
        'h207: dout <= -'sd834; // 519
        'h208: dout <=  'sd159; // 520
        'h209: dout <= -'sd236; // 521
        'h20a: dout <=  'sd7; // 522
        'h20b: dout <= -'sd378; // 523
        'h20c: dout <= -'sd1526; // 524
        'h20d: dout <= -'sd480; // 525
        'h20e: dout <= -'sd509; // 526
        'h20f: dout <= -'sd1374; // 527
        'h210: dout <=  'sd1455; // 528
        'h211: dout <= -'sd643; // 529
        'h212: dout <= -'sd1600; // 530
        'h213: dout <=  'sd307; // 531
        'h214: dout <=  'sd1583; // 532
        'h215: dout <=  'sd1288; // 533
        'h216: dout <=  'sd560; // 534
        'h217: dout <=  'sd1061; // 535
        'h218: dout <= -'sd752; // 536
        'h219: dout <= -'sd1640; // 537
        'h21a: dout <= -'sd1125; // 538
        'h21b: dout <= -'sd692; // 539
        'h21c: dout <= -'sd1014; // 540
        'h21d: dout <= -'sd148; // 541
        'h21e: dout <= -'sd1611; // 542
        'h21f: dout <= -'sd1697; // 543
        'h220: dout <= -'sd1135; // 544
        'h221: dout <= -'sd1393; // 545
        'h222: dout <=  'sd1385; // 546
        'h223: dout <=  'sd172; // 547
        'h224: dout <= -'sd1385; // 548
        'h225: dout <= -'sd325; // 549
        'h226: dout <=  'sd1707; // 550
        'h227: dout <=  'sd356; // 551
        'h228: dout <=  'sd248; // 552
        'h229: dout <= -'sd499; // 553
        'h22a: dout <= -'sd1396; // 554
        'h22b: dout <=  'sd576; // 555
        'h22c: dout <= -'sd1941; // 556
        'h22d: dout <=  'sd1314; // 557
        'h22e: dout <= -'sd2031; // 558
        'h22f: dout <=  'sd1131; // 559
        'h230: dout <= -'sd539; // 560
        'h231: dout <=  'sd837; // 561
        'h232: dout <=  'sd418; // 562
        'h233: dout <= -'sd1702; // 563
        'h234: dout <=  'sd177; // 564
        'h235: dout <= -'sd1955; // 565
        'h236: dout <= -'sd1188; // 566
        'h237: dout <= -'sd543; // 567
        'h238: dout <= -'sd984; // 568
        'h239: dout <=  'sd743; // 569
        'h23a: dout <=  'sd2235; // 570
        'h23b: dout <= -'sd657; // 571
        'h23c: dout <=  'sd1554; // 572
        'h23d: dout <= -'sd1262; // 573
        'h23e: dout <=  'sd961; // 574
        'h23f: dout <= -'sd699; // 575
        'h240: dout <=  'sd162; // 576
        'h241: dout <= -'sd1889; // 577
        'h242: dout <=  'sd1503; // 578
        'h243: dout <= -'sd1337; // 579
        'h244: dout <= -'sd168; // 580
        'h245: dout <= -'sd963; // 581
        'h246: dout <=  'sd1424; // 582
        'h247: dout <=  'sd425; // 583
        'h248: dout <=  'sd529; // 584
        'h249: dout <=  'sd1170; // 585
        'h24a: dout <= -'sd1125; // 586
        'h24b: dout <= -'sd2028; // 587
        'h24c: dout <=  'sd1508; // 588
        'h24d: dout <= -'sd847; // 589
        'h24e: dout <=  'sd1434; // 590
        'h24f: dout <=  'sd2096; // 591
        'h250: dout <=  'sd593; // 592
        'h251: dout <= -'sd1821; // 593
        'h252: dout <=  'sd1625; // 594
        'h253: dout <=  'sd613; // 595
        'h254: dout <= -'sd1167; // 596
        'h255: dout <= -'sd1341; // 597
        'h256: dout <=  'sd35; // 598
        'h257: dout <= -'sd1737; // 599
        'h258: dout <=  'sd1864; // 600
        'h259: dout <=  'sd954; // 601
        'h25a: dout <=  'sd1466; // 602
        'h25b: dout <= -'sd533; // 603
        'h25c: dout <=  'sd1943; // 604
        'h25d: dout <= -'sd1681; // 605
        'h25e: dout <=  'sd993; // 606
        'h25f: dout <= -'sd1127; // 607
        'h260: dout <= -'sd2279; // 608
        'h261: dout <= -'sd1740; // 609
        'h262: dout <= -'sd1370; // 610
        'h263: dout <=  'sd1209; // 611
        'h264: dout <= -'sd560; // 612
        'h265: dout <= -'sd82; // 613
        'h266: dout <=  'sd521; // 614
        'h267: dout <= -'sd1067; // 615
        'h268: dout <=  'sd636; // 616
        'h269: dout <=  'sd788; // 617
        'h26a: dout <=  'sd1935; // 618
        'h26b: dout <=  'sd13; // 619
        'h26c: dout <=  'sd1631; // 620
        'h26d: dout <=  'sd2147; // 621
        'h26e: dout <=  'sd1234; // 622
        'h26f: dout <= -'sd362; // 623
        'h270: dout <= -'sd1047; // 624
        'h271: dout <= -'sd1847; // 625
        'h272: dout <=  'sd1520; // 626
        'h273: dout <= -'sd1701; // 627
        'h274: dout <=  'sd273; // 628
        'h275: dout <= -'sd212; // 629
        'h276: dout <= -'sd2090; // 630
        'h277: dout <= -'sd1311; // 631
        'h278: dout <=  'sd1482; // 632
        'h279: dout <=  'sd177; // 633
        'h27a: dout <=  'sd1948; // 634
        'h27b: dout <=  'sd1873; // 635
        'h27c: dout <= -'sd1864; // 636
        'h27d: dout <=  'sd818; // 637
        'h27e: dout <= -'sd2100; // 638
        'h27f: dout <= -'sd355; // 639
        'h280: dout <= -'sd267; // 640
        'h281: dout <=  'sd2098; // 641
        'h282: dout <=  'sd438; // 642
        'h283: dout <= -'sd1423; // 643
        'h284: dout <=  'sd45; // 644
        'h285: dout <=  'sd100; // 645
        'h286: dout <= -'sd1391; // 646
        'h287: dout <= -'sd644; // 647
        'h288: dout <=  'sd1733; // 648
        'h289: dout <=  'sd2210; // 649
        'h28a: dout <=  'sd1271; // 650
        'h28b: dout <= -'sd1999; // 651
        'h28c: dout <=  'sd1863; // 652
        'h28d: dout <= -'sd191; // 653
        'h28e: dout <=  'sd1534; // 654
        'h28f: dout <= -'sd1484; // 655
        'h290: dout <= -'sd1617; // 656
        'h291: dout <=  'sd1867; // 657
        'h292: dout <= -'sd985; // 658
        'h293: dout <= -'sd2098; // 659
        'h294: dout <=  'sd5; // 660
        'h295: dout <=  'sd2252; // 661
        'h296: dout <=  'sd1540; // 662
        'h297: dout <= -'sd476; // 663
        'h298: dout <=  'sd2264; // 664
        'h299: dout <=  'sd1362; // 665
        'h29a: dout <=  'sd1570; // 666
        'h29b: dout <=  'sd671; // 667
        'h29c: dout <= -'sd485; // 668
        'h29d: dout <=  'sd1863; // 669
        'h29e: dout <= -'sd135; // 670
        'h29f: dout <=  'sd1995; // 671
        'h2a0: dout <=  'sd240; // 672
        'h2a1: dout <=  'sd1882; // 673
        'h2a2: dout <= -'sd105; // 674
        'h2a3: dout <= -'sd336; // 675
        'h2a4: dout <=  'sd407; // 676
        'h2a5: dout <= -'sd839; // 677
        'h2a6: dout <= -'sd1610; // 678
        'h2a7: dout <=  'sd410; // 679
        'h2a8: dout <=  'sd1611; // 680
        'h2a9: dout <= -'sd1020; // 681
        'h2aa: dout <=  'sd1676; // 682
        'h2ab: dout <=  'sd1318; // 683
        'h2ac: dout <=  'sd1266; // 684
        'h2ad: dout <= -'sd390; // 685
        'h2ae: dout <=  'sd2290; // 686
        'h2af: dout <=  'sd1335; // 687
        'h2b0: dout <=  'sd347; // 688
        'h2b1: dout <= -'sd1774; // 689
        'h2b2: dout <=  'sd339; // 690
        'h2b3: dout <= -'sd2229; // 691
        'h2b4: dout <=  'sd1847; // 692
        'h2b5: dout <= -'sd750; // 693
        'h2b6: dout <= -'sd604; // 694
        'h2b7: dout <=  'sd234; // 695
        'h2b8: dout <=  'sd631; // 696
        'h2b9: dout <=  'sd380; // 697
        'h2ba: dout <= -'sd69; // 698
        'h2bb: dout <=  'sd617; // 699
        'h2bc: dout <=  'sd1594; // 700
        'h2bd: dout <= -'sd247; // 701
        'h2be: dout <=  'sd0; // 702
        'h2bf: dout <=  'sd1425; // 703
        'h2c0: dout <= -'sd2280; // 704
        'h2c1: dout <= -'sd1558; // 705
        'h2c2: dout <= -'sd803; // 706
        'h2c3: dout <= -'sd1313; // 707
        'h2c4: dout <=  'sd1818; // 708
        'h2c5: dout <= -'sd1615; // 709
        'h2c6: dout <= -'sd1800; // 710
        'h2c7: dout <= -'sd839; // 711
        'h2c8: dout <=  'sd40; // 712
        'h2c9: dout <=  'sd1476; // 713
        'h2ca: dout <=  'sd2276; // 714
        'h2cb: dout <=  'sd1615; // 715
        'h2cc: dout <=  'sd500; // 716
        'h2cd: dout <= -'sd2123; // 717
        'h2ce: dout <= -'sd2004; // 718
        'h2cf: dout <=  'sd600; // 719
        'h2d0: dout <=  'sd1469; // 720
        'h2d1: dout <= -'sd1077; // 721
        'h2d2: dout <=  'sd2154; // 722
        'h2d3: dout <=  'sd231; // 723
        'h2d4: dout <=  'sd339; // 724
        'h2d5: dout <=  'sd545; // 725
        'h2d6: dout <= -'sd1952; // 726
        'h2d7: dout <= -'sd1513; // 727
        'h2d8: dout <=  'sd2003; // 728
        'h2d9: dout <= -'sd1068; // 729
        'h2da: dout <= -'sd1913; // 730
        'h2db: dout <= -'sd999; // 731
        'h2dc: dout <=  'sd1038; // 732
        'h2dd: dout <= -'sd1089; // 733
        'h2de: dout <= -'sd1329; // 734
        'h2df: dout <= -'sd1023; // 735
        'h2e0: dout <= -'sd90; // 736
        'h2e1: dout <=  'sd1091; // 737
        'h2e2: dout <= -'sd912; // 738
        'h2e3: dout <=  'sd1715; // 739
        'h2e4: dout <=  'sd2185; // 740
        'h2e5: dout <=  'sd1478; // 741
        'h2e6: dout <= -'sd1951; // 742
        'h2e7: dout <= -'sd847; // 743
        'h2e8: dout <=  'sd1955; // 744
        'h2e9: dout <=  'sd1650; // 745
        'h2ea: dout <= -'sd1684; // 746
        'h2eb: dout <= -'sd265; // 747
        'h2ec: dout <= -'sd625; // 748
        'h2ed: dout <=  'sd1136; // 749
        'h2ee: dout <= -'sd2164; // 750
        'h2ef: dout <= -'sd847; // 751
        'h2f0: dout <=  'sd1147; // 752
        'h2f1: dout <=  'sd1776; // 753
        'h2f2: dout <= -'sd2109; // 754
        'h2f3: dout <=  'sd406; // 755
        'h2f4: dout <=  'sd751; // 756
        'h2f5: dout <=  'sd1712; // 757
        'h2f6: dout <= -'sd346; // 758
        'h2f7: dout <=  'sd2172; // 759
        'h2f8: dout <= -'sd1389; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module h_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <=  'sd1418; // 0
        'h001: dout <=  'sd2023; // 1
        'h002: dout <=  'sd178; // 2
        'h003: dout <= -'sd1610; // 3
        'h004: dout <=  'sd494; // 4
        'h005: dout <= -'sd1848; // 5
        'h006: dout <=  'sd2039; // 6
        'h007: dout <=  'sd342; // 7
        'h008: dout <=  'sd2165; // 8
        'h009: dout <= -'sd390; // 9
        'h00a: dout <=  'sd1777; // 10
        'h00b: dout <=  'sd2068; // 11
        'h00c: dout <=  'sd1687; // 12
        'h00d: dout <=  'sd2154; // 13
        'h00e: dout <=  'sd1503; // 14
        'h00f: dout <=  'sd1076; // 15
        'h010: dout <= -'sd1472; // 16
        'h011: dout <=  'sd935; // 17
        'h012: dout <=  'sd617; // 18
        'h013: dout <= -'sd1462; // 19
        'h014: dout <=  'sd2171; // 20
        'h015: dout <= -'sd1720; // 21
        'h016: dout <= -'sd1254; // 22
        'h017: dout <=  'sd2007; // 23
        'h018: dout <=  'sd817; // 24
        'h019: dout <= -'sd32; // 25
        'h01a: dout <= -'sd604; // 26
        'h01b: dout <=  'sd2133; // 27
        'h01c: dout <= -'sd1366; // 28
        'h01d: dout <= -'sd1098; // 29
        'h01e: dout <= -'sd382; // 30
        'h01f: dout <= -'sd2072; // 31
        'h020: dout <=  'sd416; // 32
        'h021: dout <=  'sd217; // 33
        'h022: dout <= -'sd1153; // 34
        'h023: dout <= -'sd352; // 35
        'h024: dout <= -'sd1261; // 36
        'h025: dout <= -'sd1586; // 37
        'h026: dout <=  'sd255; // 38
        'h027: dout <= -'sd690; // 39
        'h028: dout <=  'sd1783; // 40
        'h029: dout <= -'sd318; // 41
        'h02a: dout <= -'sd1741; // 42
        'h02b: dout <= -'sd906; // 43
        'h02c: dout <=  'sd15; // 44
        'h02d: dout <= -'sd2041; // 45
        'h02e: dout <=  'sd1736; // 46
        'h02f: dout <= -'sd1396; // 47
        'h030: dout <= -'sd1433; // 48
        'h031: dout <=  'sd490; // 49
        'h032: dout <= -'sd622; // 50
        'h033: dout <= -'sd1928; // 51
        'h034: dout <= -'sd640; // 52
        'h035: dout <= -'sd1030; // 53
        'h036: dout <=  'sd722; // 54
        'h037: dout <= -'sd860; // 55
        'h038: dout <=  'sd1373; // 56
        'h039: dout <=  'sd1103; // 57
        'h03a: dout <= -'sd582; // 58
        'h03b: dout <= -'sd918; // 59
        'h03c: dout <=  'sd802; // 60
        'h03d: dout <=  'sd1762; // 61
        'h03e: dout <=  'sd1084; // 62
        'h03f: dout <=  'sd1652; // 63
        'h040: dout <=  'sd248; // 64
        'h041: dout <=  'sd277; // 65
        'h042: dout <=  'sd944; // 66
        'h043: dout <= -'sd540; // 67
        'h044: dout <= -'sd81; // 68
        'h045: dout <= -'sd1789; // 69
        'h046: dout <= -'sd687; // 70
        'h047: dout <=  'sd2052; // 71
        'h048: dout <= -'sd598; // 72
        'h049: dout <=  'sd1420; // 73
        'h04a: dout <=  'sd1964; // 74
        'h04b: dout <=  'sd389; // 75
        'h04c: dout <= -'sd358; // 76
        'h04d: dout <=  'sd1511; // 77
        'h04e: dout <= -'sd869; // 78
        'h04f: dout <=  'sd1554; // 79
        'h050: dout <= -'sd843; // 80
        'h051: dout <= -'sd64; // 81
        'h052: dout <=  'sd225; // 82
        'h053: dout <= -'sd1288; // 83
        'h054: dout <= -'sd1300; // 84
        'h055: dout <= -'sd2063; // 85
        'h056: dout <= -'sd1235; // 86
        'h057: dout <=  'sd1683; // 87
        'h058: dout <= -'sd1750; // 88
        'h059: dout <=  'sd34; // 89
        'h05a: dout <=  'sd25; // 90
        'h05b: dout <=  'sd1439; // 91
        'h05c: dout <= -'sd1359; // 92
        'h05d: dout <= -'sd1410; // 93
        'h05e: dout <=  'sd314; // 94
        'h05f: dout <= -'sd464; // 95
        'h060: dout <=  'sd1101; // 96
        'h061: dout <=  'sd1031; // 97
        'h062: dout <= -'sd1221; // 98
        'h063: dout <=  'sd197; // 99
        'h064: dout <= -'sd1950; // 100
        'h065: dout <=  'sd506; // 101
        'h066: dout <=  'sd2266; // 102
        'h067: dout <=  'sd1016; // 103
        'h068: dout <=  'sd1917; // 104
        'h069: dout <= -'sd1219; // 105
        'h06a: dout <=  'sd192; // 106
        'h06b: dout <=  'sd1132; // 107
        'h06c: dout <= -'sd1118; // 108
        'h06d: dout <=  'sd1327; // 109
        'h06e: dout <=  'sd1866; // 110
        'h06f: dout <= -'sd1110; // 111
        'h070: dout <=  'sd1924; // 112
        'h071: dout <= -'sd179; // 113
        'h072: dout <= -'sd776; // 114
        'h073: dout <=  'sd4; // 115
        'h074: dout <=  'sd2061; // 116
        'h075: dout <=  'sd2129; // 117
        'h076: dout <= -'sd2171; // 118
        'h077: dout <=  'sd974; // 119
        'h078: dout <=  'sd235; // 120
        'h079: dout <= -'sd64; // 121
        'h07a: dout <=  'sd672; // 122
        'h07b: dout <= -'sd1481; // 123
        'h07c: dout <= -'sd151; // 124
        'h07d: dout <=  'sd866; // 125
        'h07e: dout <= -'sd1616; // 126
        'h07f: dout <= -'sd1128; // 127
        'h080: dout <= -'sd770; // 128
        'h081: dout <=  'sd196; // 129
        'h082: dout <= -'sd2187; // 130
        'h083: dout <= -'sd1110; // 131
        'h084: dout <=  'sd1513; // 132
        'h085: dout <=  'sd2096; // 133
        'h086: dout <=  'sd695; // 134
        'h087: dout <=  'sd841; // 135
        'h088: dout <=  'sd648; // 136
        'h089: dout <=  'sd192; // 137
        'h08a: dout <=  'sd1301; // 138
        'h08b: dout <= -'sd1912; // 139
        'h08c: dout <= -'sd1231; // 140
        'h08d: dout <= -'sd2170; // 141
        'h08e: dout <=  'sd179; // 142
        'h08f: dout <= -'sd87; // 143
        'h090: dout <=  'sd2057; // 144
        'h091: dout <= -'sd2222; // 145
        'h092: dout <=  'sd164; // 146
        'h093: dout <= -'sd716; // 147
        'h094: dout <= -'sd1922; // 148
        'h095: dout <=  'sd372; // 149
        'h096: dout <=  'sd250; // 150
        'h097: dout <= -'sd483; // 151
        'h098: dout <=  'sd779; // 152
        'h099: dout <= -'sd1379; // 153
        'h09a: dout <= -'sd538; // 154
        'h09b: dout <=  'sd91; // 155
        'h09c: dout <= -'sd1042; // 156
        'h09d: dout <= -'sd1592; // 157
        'h09e: dout <=  'sd1256; // 158
        'h09f: dout <= -'sd903; // 159
        'h0a0: dout <= -'sd433; // 160
        'h0a1: dout <= -'sd1236; // 161
        'h0a2: dout <= -'sd1281; // 162
        'h0a3: dout <=  'sd2249; // 163
        'h0a4: dout <=  'sd241; // 164
        'h0a5: dout <=  'sd1776; // 165
        'h0a6: dout <=  'sd1503; // 166
        'h0a7: dout <= -'sd1425; // 167
        'h0a8: dout <= -'sd642; // 168
        'h0a9: dout <=  'sd308; // 169
        'h0aa: dout <=  'sd123; // 170
        'h0ab: dout <=  'sd191; // 171
        'h0ac: dout <= -'sd622; // 172
        'h0ad: dout <= -'sd855; // 173
        'h0ae: dout <=  'sd143; // 174
        'h0af: dout <=  'sd1849; // 175
        'h0b0: dout <=  'sd64; // 176
        'h0b1: dout <= -'sd958; // 177
        'h0b2: dout <=  'sd251; // 178
        'h0b3: dout <=  'sd452; // 179
        'h0b4: dout <=  'sd1351; // 180
        'h0b5: dout <= -'sd2075; // 181
        'h0b6: dout <= -'sd1264; // 182
        'h0b7: dout <=  'sd1122; // 183
        'h0b8: dout <=  'sd937; // 184
        'h0b9: dout <= -'sd1350; // 185
        'h0ba: dout <= -'sd93; // 186
        'h0bb: dout <=  'sd1002; // 187
        'h0bc: dout <= -'sd646; // 188
        'h0bd: dout <= -'sd1811; // 189
        'h0be: dout <= -'sd1388; // 190
        'h0bf: dout <=  'sd612; // 191
        'h0c0: dout <= -'sd2080; // 192
        'h0c1: dout <= -'sd396; // 193
        'h0c2: dout <= -'sd1206; // 194
        'h0c3: dout <=  'sd1380; // 195
        'h0c4: dout <= -'sd1680; // 196
        'h0c5: dout <= -'sd819; // 197
        'h0c6: dout <= -'sd1827; // 198
        'h0c7: dout <=  'sd2250; // 199
        'h0c8: dout <=  'sd1599; // 200
        'h0c9: dout <= -'sd755; // 201
        'h0ca: dout <=  'sd640; // 202
        'h0cb: dout <= -'sd547; // 203
        'h0cc: dout <= -'sd1881; // 204
        'h0cd: dout <=  'sd1534; // 205
        'h0ce: dout <= -'sd2052; // 206
        'h0cf: dout <=  'sd912; // 207
        'h0d0: dout <=  'sd2232; // 208
        'h0d1: dout <= -'sd169; // 209
        'h0d2: dout <=  'sd1418; // 210
        'h0d3: dout <= -'sd416; // 211
        'h0d4: dout <=  'sd1979; // 212
        'h0d5: dout <= -'sd54; // 213
        'h0d6: dout <=  'sd431; // 214
        'h0d7: dout <= -'sd2220; // 215
        'h0d8: dout <=  'sd1764; // 216
        'h0d9: dout <=  'sd1666; // 217
        'h0da: dout <= -'sd771; // 218
        'h0db: dout <= -'sd1673; // 219
        'h0dc: dout <= -'sd1316; // 220
        'h0dd: dout <= -'sd1065; // 221
        'h0de: dout <=  'sd821; // 222
        'h0df: dout <=  'sd143; // 223
        'h0e0: dout <= -'sd1189; // 224
        'h0e1: dout <=  'sd643; // 225
        'h0e2: dout <=  'sd1157; // 226
        'h0e3: dout <=  'sd1877; // 227
        'h0e4: dout <=  'sd853; // 228
        'h0e5: dout <=  'sd1954; // 229
        'h0e6: dout <=  'sd723; // 230
        'h0e7: dout <=  'sd1956; // 231
        'h0e8: dout <=  'sd1094; // 232
        'h0e9: dout <= -'sd83; // 233
        'h0ea: dout <= -'sd472; // 234
        'h0eb: dout <= -'sd1354; // 235
        'h0ec: dout <= -'sd586; // 236
        'h0ed: dout <= -'sd1209; // 237
        'h0ee: dout <= -'sd1377; // 238
        'h0ef: dout <=  'sd48; // 239
        'h0f0: dout <=  'sd1161; // 240
        'h0f1: dout <=  'sd1307; // 241
        'h0f2: dout <=  'sd1668; // 242
        'h0f3: dout <=  'sd438; // 243
        'h0f4: dout <=  'sd1704; // 244
        'h0f5: dout <=  'sd670; // 245
        'h0f6: dout <= -'sd1328; // 246
        'h0f7: dout <=  'sd541; // 247
        'h0f8: dout <=  'sd914; // 248
        'h0f9: dout <= -'sd1935; // 249
        'h0fa: dout <=  'sd2032; // 250
        'h0fb: dout <= -'sd2068; // 251
        'h0fc: dout <=  'sd1927; // 252
        'h0fd: dout <= -'sd1810; // 253
        'h0fe: dout <= -'sd1331; // 254
        'h0ff: dout <= -'sd1867; // 255
        'h100: dout <=  'sd750; // 256
        'h101: dout <= -'sd361; // 257
        'h102: dout <= -'sd565; // 258
        'h103: dout <= -'sd1077; // 259
        'h104: dout <=  'sd1875; // 260
        'h105: dout <=  'sd947; // 261
        'h106: dout <=  'sd850; // 262
        'h107: dout <=  'sd131; // 263
        'h108: dout <=  'sd1505; // 264
        'h109: dout <=  'sd1463; // 265
        'h10a: dout <=  'sd907; // 266
        'h10b: dout <=  'sd295; // 267
        'h10c: dout <= -'sd1484; // 268
        'h10d: dout <=  'sd1511; // 269
        'h10e: dout <=  'sd808; // 270
        'h10f: dout <= -'sd1801; // 271
        'h110: dout <=  'sd2034; // 272
        'h111: dout <=  'sd110; // 273
        'h112: dout <= -'sd2106; // 274
        'h113: dout <= -'sd910; // 275
        'h114: dout <= -'sd1056; // 276
        'h115: dout <= -'sd1311; // 277
        'h116: dout <= -'sd1733; // 278
        'h117: dout <= -'sd1119; // 279
        'h118: dout <= -'sd11; // 280
        'h119: dout <= -'sd1562; // 281
        'h11a: dout <= -'sd895; // 282
        'h11b: dout <= -'sd207; // 283
        'h11c: dout <=  'sd1606; // 284
        'h11d: dout <= -'sd635; // 285
        'h11e: dout <=  'sd163; // 286
        'h11f: dout <=  'sd2076; // 287
        'h120: dout <= -'sd2082; // 288
        'h121: dout <= -'sd1813; // 289
        'h122: dout <= -'sd445; // 290
        'h123: dout <=  'sd1871; // 291
        'h124: dout <=  'sd2243; // 292
        'h125: dout <=  'sd650; // 293
        'h126: dout <= -'sd172; // 294
        'h127: dout <=  'sd1419; // 295
        'h128: dout <= -'sd1231; // 296
        'h129: dout <= -'sd2170; // 297
        'h12a: dout <=  'sd123; // 298
        'h12b: dout <= -'sd405; // 299
        'h12c: dout <=  'sd1834; // 300
        'h12d: dout <=  'sd580; // 301
        'h12e: dout <= -'sd1272; // 302
        'h12f: dout <= -'sd1299; // 303
        'h130: dout <=  'sd1781; // 304
        'h131: dout <=  'sd1006; // 305
        'h132: dout <= -'sd319; // 306
        'h133: dout <=  'sd1402; // 307
        'h134: dout <= -'sd1695; // 308
        'h135: dout <=  'sd1266; // 309
        'h136: dout <=  'sd1026; // 310
        'h137: dout <= -'sd251; // 311
        'h138: dout <= -'sd869; // 312
        'h139: dout <=  'sd1314; // 313
        'h13a: dout <=  'sd1525; // 314
        'h13b: dout <= -'sd1239; // 315
        'h13c: dout <= -'sd558; // 316
        'h13d: dout <=  'sd1773; // 317
        'h13e: dout <= -'sd518; // 318
        'h13f: dout <=  'sd459; // 319
        'h140: dout <= -'sd1964; // 320
        'h141: dout <=  'sd134; // 321
        'h142: dout <=  'sd154; // 322
        'h143: dout <= -'sd1988; // 323
        'h144: dout <= -'sd1733; // 324
        'h145: dout <=  'sd732; // 325
        'h146: dout <=  'sd1017; // 326
        'h147: dout <=  'sd1960; // 327
        'h148: dout <= -'sd1191; // 328
        'h149: dout <=  'sd52; // 329
        'h14a: dout <= -'sd1065; // 330
        'h14b: dout <= -'sd714; // 331
        'h14c: dout <= -'sd981; // 332
        'h14d: dout <=  'sd1389; // 333
        'h14e: dout <=  'sd1530; // 334
        'h14f: dout <=  'sd738; // 335
        'h150: dout <= -'sd8; // 336
        'h151: dout <= -'sd1873; // 337
        'h152: dout <= -'sd1380; // 338
        'h153: dout <=  'sd860; // 339
        'h154: dout <= -'sd1548; // 340
        'h155: dout <=  'sd109; // 341
        'h156: dout <=  'sd1073; // 342
        'h157: dout <=  'sd1789; // 343
        'h158: dout <= -'sd427; // 344
        'h159: dout <=  'sd242; // 345
        'h15a: dout <=  'sd271; // 346
        'h15b: dout <=  'sd2274; // 347
        'h15c: dout <=  'sd1264; // 348
        'h15d: dout <= -'sd2128; // 349
        'h15e: dout <= -'sd434; // 350
        'h15f: dout <= -'sd1294; // 351
        'h160: dout <=  'sd1419; // 352
        'h161: dout <= -'sd1421; // 353
        'h162: dout <=  'sd1711; // 354
        'h163: dout <= -'sd1381; // 355
        'h164: dout <= -'sd119; // 356
        'h165: dout <= -'sd1250; // 357
        'h166: dout <= -'sd1664; // 358
        'h167: dout <= -'sd844; // 359
        'h168: dout <=  'sd1309; // 360
        'h169: dout <=  'sd1745; // 361
        'h16a: dout <= -'sd1066; // 362
        'h16b: dout <= -'sd1878; // 363
        'h16c: dout <=  'sd436; // 364
        'h16d: dout <= -'sd1384; // 365
        'h16e: dout <= -'sd532; // 366
        'h16f: dout <=  'sd1084; // 367
        'h170: dout <=  'sd655; // 368
        'h171: dout <= -'sd796; // 369
        'h172: dout <=  'sd600; // 370
        'h173: dout <= -'sd2135; // 371
        'h174: dout <= -'sd138; // 372
        'h175: dout <= -'sd1344; // 373
        'h176: dout <=  'sd295; // 374
        'h177: dout <=  'sd1716; // 375
        'h178: dout <= -'sd513; // 376
        'h179: dout <= -'sd511; // 377
        'h17a: dout <= -'sd2088; // 378
        'h17b: dout <= -'sd776; // 379
        'h17c: dout <=  'sd762; // 380
        'h17d: dout <= -'sd487; // 381
        'h17e: dout <=  'sd556; // 382
        'h17f: dout <=  'sd1399; // 383
        'h180: dout <=  'sd155; // 384
        'h181: dout <= -'sd714; // 385
        'h182: dout <= -'sd794; // 386
        'h183: dout <= -'sd893; // 387
        'h184: dout <= -'sd1341; // 388
        'h185: dout <= -'sd1068; // 389
        'h186: dout <=  'sd2053; // 390
        'h187: dout <= -'sd1617; // 391
        'h188: dout <=  'sd365; // 392
        'h189: dout <=  'sd848; // 393
        'h18a: dout <=  'sd321; // 394
        'h18b: dout <=  'sd1691; // 395
        'h18c: dout <=  'sd979; // 396
        'h18d: dout <= -'sd1499; // 397
        'h18e: dout <=  'sd1203; // 398
        'h18f: dout <=  'sd1720; // 399
        'h190: dout <= -'sd548; // 400
        'h191: dout <=  'sd1391; // 401
        'h192: dout <= -'sd1629; // 402
        'h193: dout <= -'sd195; // 403
        'h194: dout <=  'sd879; // 404
        'h195: dout <=  'sd1952; // 405
        'h196: dout <=  'sd1588; // 406
        'h197: dout <=  'sd1318; // 407
        'h198: dout <=  'sd103; // 408
        'h199: dout <=  'sd2257; // 409
        'h19a: dout <=  'sd948; // 410
        'h19b: dout <=  'sd1354; // 411
        'h19c: dout <=  'sd247; // 412
        'h19d: dout <= -'sd1636; // 413
        'h19e: dout <=  'sd1114; // 414
        'h19f: dout <= -'sd196; // 415
        'h1a0: dout <=  'sd1505; // 416
        'h1a1: dout <= -'sd1737; // 417
        'h1a2: dout <=  'sd980; // 418
        'h1a3: dout <=  'sd1577; // 419
        'h1a4: dout <= -'sd398; // 420
        'h1a5: dout <=  'sd542; // 421
        'h1a6: dout <=  'sd613; // 422
        'h1a7: dout <=  'sd303; // 423
        'h1a8: dout <=  'sd2242; // 424
        'h1a9: dout <= -'sd2233; // 425
        'h1aa: dout <=  'sd2067; // 426
        'h1ab: dout <=  'sd786; // 427
        'h1ac: dout <= -'sd1077; // 428
        'h1ad: dout <=  'sd1698; // 429
        'h1ae: dout <=  'sd556; // 430
        'h1af: dout <=  'sd2023; // 431
        'h1b0: dout <=  'sd1306; // 432
        'h1b1: dout <=  'sd1175; // 433
        'h1b2: dout <=  'sd1968; // 434
        'h1b3: dout <=  'sd116; // 435
        'h1b4: dout <=  'sd169; // 436
        'h1b5: dout <=  'sd676; // 437
        'h1b6: dout <=  'sd482; // 438
        'h1b7: dout <= -'sd517; // 439
        'h1b8: dout <= -'sd618; // 440
        'h1b9: dout <= -'sd1147; // 441
        'h1ba: dout <=  'sd1296; // 442
        'h1bb: dout <= -'sd471; // 443
        'h1bc: dout <= -'sd446; // 444
        'h1bd: dout <=  'sd492; // 445
        'h1be: dout <=  'sd2209; // 446
        'h1bf: dout <=  'sd962; // 447
        'h1c0: dout <= -'sd2021; // 448
        'h1c1: dout <= -'sd787; // 449
        'h1c2: dout <= -'sd1023; // 450
        'h1c3: dout <=  'sd1228; // 451
        'h1c4: dout <=  'sd1505; // 452
        'h1c5: dout <= -'sd1497; // 453
        'h1c6: dout <=  'sd1477; // 454
        'h1c7: dout <=  'sd710; // 455
        'h1c8: dout <= -'sd528; // 456
        'h1c9: dout <=  'sd443; // 457
        'h1ca: dout <=  'sd1797; // 458
        'h1cb: dout <=  'sd524; // 459
        'h1cc: dout <= -'sd1758; // 460
        'h1cd: dout <= -'sd1779; // 461
        'h1ce: dout <= -'sd764; // 462
        'h1cf: dout <=  'sd1727; // 463
        'h1d0: dout <= -'sd1133; // 464
        'h1d1: dout <= -'sd390; // 465
        'h1d2: dout <=  'sd1395; // 466
        'h1d3: dout <=  'sd224; // 467
        'h1d4: dout <= -'sd1717; // 468
        'h1d5: dout <=  'sd2106; // 469
        'h1d6: dout <= -'sd52; // 470
        'h1d7: dout <= -'sd1533; // 471
        'h1d8: dout <=  'sd776; // 472
        'h1d9: dout <= -'sd1011; // 473
        'h1da: dout <= -'sd225; // 474
        'h1db: dout <=  'sd593; // 475
        'h1dc: dout <= -'sd897; // 476
        'h1dd: dout <=  'sd1934; // 477
        'h1de: dout <= -'sd1774; // 478
        'h1df: dout <=  'sd1759; // 479
        'h1e0: dout <= -'sd857; // 480
        'h1e1: dout <=  'sd1096; // 481
        'h1e2: dout <= -'sd1352; // 482
        'h1e3: dout <=  'sd1247; // 483
        'h1e4: dout <=  'sd1642; // 484
        'h1e5: dout <=  'sd1723; // 485
        'h1e6: dout <=  'sd1388; // 486
        'h1e7: dout <= -'sd562; // 487
        'h1e8: dout <= -'sd1516; // 488
        'h1e9: dout <=  'sd1775; // 489
        'h1ea: dout <=  'sd2196; // 490
        'h1eb: dout <=  'sd322; // 491
        'h1ec: dout <=  'sd2164; // 492
        'h1ed: dout <= -'sd1045; // 493
        'h1ee: dout <=  'sd465; // 494
        'h1ef: dout <=  'sd1361; // 495
        'h1f0: dout <=  'sd90; // 496
        'h1f1: dout <=  'sd1885; // 497
        'h1f2: dout <=  'sd590; // 498
        'h1f3: dout <=  'sd486; // 499
        'h1f4: dout <= -'sd1477; // 500
        'h1f5: dout <=  'sd661; // 501
        'h1f6: dout <= -'sd129; // 502
        'h1f7: dout <=  'sd1487; // 503
        'h1f8: dout <=  'sd655; // 504
        'h1f9: dout <= -'sd1386; // 505
        'h1fa: dout <=  'sd1572; // 506
        'h1fb: dout <= -'sd984; // 507
        'h1fc: dout <= -'sd1158; // 508
        'h1fd: dout <=  'sd1038; // 509
        'h1fe: dout <= -'sd690; // 510
        'h1ff: dout <=  'sd1614; // 511
        'h200: dout <=  'sd2172; // 512
        'h201: dout <=  'sd928; // 513
        'h202: dout <= -'sd1616; // 514
        'h203: dout <=  'sd1978; // 515
        'h204: dout <= -'sd1026; // 516
        'h205: dout <= -'sd739; // 517
        'h206: dout <= -'sd1881; // 518
        'h207: dout <=  'sd2124; // 519
        'h208: dout <=  'sd1608; // 520
        'h209: dout <=  'sd2254; // 521
        'h20a: dout <=  'sd943; // 522
        'h20b: dout <=  'sd643; // 523
        'h20c: dout <=  'sd795; // 524
        'h20d: dout <= -'sd1451; // 525
        'h20e: dout <=  'sd1275; // 526
        'h20f: dout <= -'sd689; // 527
        'h210: dout <= -'sd835; // 528
        'h211: dout <=  'sd2175; // 529
        'h212: dout <= -'sd1342; // 530
        'h213: dout <=  'sd762; // 531
        'h214: dout <= -'sd1965; // 532
        'h215: dout <=  'sd1366; // 533
        'h216: dout <=  'sd2065; // 534
        'h217: dout <=  'sd836; // 535
        'h218: dout <= -'sd237; // 536
        'h219: dout <=  'sd1353; // 537
        'h21a: dout <= -'sd298; // 538
        'h21b: dout <=  'sd453; // 539
        'h21c: dout <= -'sd1631; // 540
        'h21d: dout <=  'sd967; // 541
        'h21e: dout <= -'sd788; // 542
        'h21f: dout <=  'sd550; // 543
        'h220: dout <=  'sd424; // 544
        'h221: dout <=  'sd80; // 545
        'h222: dout <= -'sd1818; // 546
        'h223: dout <= -'sd1504; // 547
        'h224: dout <=  'sd143; // 548
        'h225: dout <= -'sd1751; // 549
        'h226: dout <=  'sd495; // 550
        'h227: dout <= -'sd1197; // 551
        'h228: dout <= -'sd1700; // 552
        'h229: dout <= -'sd1510; // 553
        'h22a: dout <=  'sd1960; // 554
        'h22b: dout <= -'sd1491; // 555
        'h22c: dout <=  'sd686; // 556
        'h22d: dout <= -'sd2156; // 557
        'h22e: dout <=  'sd1773; // 558
        'h22f: dout <=  'sd1006; // 559
        'h230: dout <= -'sd435; // 560
        'h231: dout <= -'sd155; // 561
        'h232: dout <=  'sd412; // 562
        'h233: dout <=  'sd1825; // 563
        'h234: dout <=  'sd1319; // 564
        'h235: dout <=  'sd743; // 565
        'h236: dout <= -'sd1246; // 566
        'h237: dout <= -'sd2254; // 567
        'h238: dout <=  'sd686; // 568
        'h239: dout <= -'sd1366; // 569
        'h23a: dout <= -'sd1284; // 570
        'h23b: dout <= -'sd1926; // 571
        'h23c: dout <= -'sd1680; // 572
        'h23d: dout <= -'sd655; // 573
        'h23e: dout <=  'sd565; // 574
        'h23f: dout <= -'sd223; // 575
        'h240: dout <=  'sd2264; // 576
        'h241: dout <=  'sd512; // 577
        'h242: dout <=  'sd997; // 578
        'h243: dout <= -'sd1370; // 579
        'h244: dout <= -'sd202; // 580
        'h245: dout <= -'sd2125; // 581
        'h246: dout <=  'sd433; // 582
        'h247: dout <=  'sd593; // 583
        'h248: dout <= -'sd521; // 584
        'h249: dout <= -'sd1484; // 585
        'h24a: dout <=  'sd588; // 586
        'h24b: dout <=  'sd859; // 587
        'h24c: dout <= -'sd1621; // 588
        'h24d: dout <=  'sd1523; // 589
        'h24e: dout <=  'sd813; // 590
        'h24f: dout <=  'sd1322; // 591
        'h250: dout <= -'sd1610; // 592
        'h251: dout <= -'sd2013; // 593
        'h252: dout <=  'sd1341; // 594
        'h253: dout <=  'sd215; // 595
        'h254: dout <=  'sd939; // 596
        'h255: dout <= -'sd2289; // 597
        'h256: dout <= -'sd1136; // 598
        'h257: dout <= -'sd39; // 599
        'h258: dout <= -'sd1525; // 600
        'h259: dout <=  'sd1519; // 601
        'h25a: dout <=  'sd2080; // 602
        'h25b: dout <=  'sd1080; // 603
        'h25c: dout <= -'sd610; // 604
        'h25d: dout <=  'sd2038; // 605
        'h25e: dout <= -'sd1303; // 606
        'h25f: dout <=  'sd2102; // 607
        'h260: dout <=  'sd667; // 608
        'h261: dout <=  'sd1764; // 609
        'h262: dout <=  'sd1106; // 610
        'h263: dout <= -'sd287; // 611
        'h264: dout <=  'sd2216; // 612
        'h265: dout <=  'sd1395; // 613
        'h266: dout <=  'sd1252; // 614
        'h267: dout <=  'sd668; // 615
        'h268: dout <= -'sd77; // 616
        'h269: dout <= -'sd1626; // 617
        'h26a: dout <= -'sd1132; // 618
        'h26b: dout <= -'sd466; // 619
        'h26c: dout <=  'sd1337; // 620
        'h26d: dout <= -'sd1711; // 621
        'h26e: dout <= -'sd460; // 622
        'h26f: dout <=  'sd1846; // 623
        'h270: dout <=  'sd1903; // 624
        'h271: dout <=  'sd1218; // 625
        'h272: dout <=  'sd1084; // 626
        'h273: dout <=  'sd285; // 627
        'h274: dout <=  'sd1877; // 628
        'h275: dout <=  'sd1739; // 629
        'h276: dout <=  'sd736; // 630
        'h277: dout <= -'sd598; // 631
        'h278: dout <= -'sd10; // 632
        'h279: dout <=  'sd1272; // 633
        'h27a: dout <= -'sd1636; // 634
        'h27b: dout <=  'sd1271; // 635
        'h27c: dout <=  'sd728; // 636
        'h27d: dout <=  'sd69; // 637
        'h27e: dout <=  'sd525; // 638
        'h27f: dout <=  'sd1093; // 639
        'h280: dout <= -'sd2231; // 640
        'h281: dout <=  'sd1366; // 641
        'h282: dout <= -'sd272; // 642
        'h283: dout <= -'sd1877; // 643
        'h284: dout <=  'sd477; // 644
        'h285: dout <= -'sd903; // 645
        'h286: dout <= -'sd774; // 646
        'h287: dout <=  'sd2217; // 647
        'h288: dout <=  'sd332; // 648
        'h289: dout <= -'sd1700; // 649
        'h28a: dout <= -'sd724; // 650
        'h28b: dout <= -'sd74; // 651
        'h28c: dout <= -'sd1682; // 652
        'h28d: dout <= -'sd1222; // 653
        'h28e: dout <= -'sd850; // 654
        'h28f: dout <= -'sd1128; // 655
        'h290: dout <=  'sd895; // 656
        'h291: dout <=  'sd98; // 657
        'h292: dout <= -'sd2135; // 658
        'h293: dout <= -'sd2160; // 659
        'h294: dout <= -'sd1319; // 660
        'h295: dout <=  'sd978; // 661
        'h296: dout <= -'sd2067; // 662
        'h297: dout <=  'sd507; // 663
        'h298: dout <=  'sd398; // 664
        'h299: dout <=  'sd316; // 665
        'h29a: dout <=  'sd267; // 666
        'h29b: dout <=  'sd1696; // 667
        'h29c: dout <= -'sd278; // 668
        'h29d: dout <=  'sd1522; // 669
        'h29e: dout <=  'sd1579; // 670
        'h29f: dout <= -'sd1984; // 671
        'h2a0: dout <=  'sd8; // 672
        'h2a1: dout <= -'sd427; // 673
        'h2a2: dout <=  'sd64; // 674
        'h2a3: dout <=  'sd1607; // 675
        'h2a4: dout <=  'sd949; // 676
        'h2a5: dout <=  'sd716; // 677
        'h2a6: dout <= -'sd2292; // 678
        'h2a7: dout <= -'sd1921; // 679
        'h2a8: dout <=  'sd1459; // 680
        'h2a9: dout <= -'sd2233; // 681
        'h2aa: dout <=  'sd1163; // 682
        'h2ab: dout <=  'sd647; // 683
        'h2ac: dout <=  'sd1984; // 684
        'h2ad: dout <= -'sd917; // 685
        'h2ae: dout <=  'sd643; // 686
        'h2af: dout <= -'sd1007; // 687
        'h2b0: dout <=  'sd1582; // 688
        'h2b1: dout <= -'sd1968; // 689
        'h2b2: dout <= -'sd1148; // 690
        'h2b3: dout <=  'sd1375; // 691
        'h2b4: dout <= -'sd1943; // 692
        'h2b5: dout <= -'sd367; // 693
        'h2b6: dout <=  'sd1930; // 694
        'h2b7: dout <=  'sd926; // 695
        'h2b8: dout <=  'sd263; // 696
        'h2b9: dout <= -'sd1357; // 697
        'h2ba: dout <= -'sd1642; // 698
        'h2bb: dout <= -'sd1223; // 699
        'h2bc: dout <=  'sd1048; // 700
        'h2bd: dout <= -'sd2084; // 701
        'h2be: dout <=  'sd177; // 702
        'h2bf: dout <= -'sd1350; // 703
        'h2c0: dout <=  'sd2130; // 704
        'h2c1: dout <=  'sd480; // 705
        'h2c2: dout <=  'sd734; // 706
        'h2c3: dout <=  'sd421; // 707
        'h2c4: dout <= -'sd1536; // 708
        'h2c5: dout <=  'sd1757; // 709
        'h2c6: dout <=  'sd303; // 710
        'h2c7: dout <= -'sd1939; // 711
        'h2c8: dout <=  'sd468; // 712
        'h2c9: dout <=  'sd973; // 713
        'h2ca: dout <=  'sd230; // 714
        'h2cb: dout <=  'sd594; // 715
        'h2cc: dout <=  'sd432; // 716
        'h2cd: dout <=  'sd577; // 717
        'h2ce: dout <=  'sd758; // 718
        'h2cf: dout <=  'sd2115; // 719
        'h2d0: dout <=  'sd268; // 720
        'h2d1: dout <= -'sd1340; // 721
        'h2d2: dout <=  'sd309; // 722
        'h2d3: dout <=  'sd1291; // 723
        'h2d4: dout <=  'sd1397; // 724
        'h2d5: dout <= -'sd1920; // 725
        'h2d6: dout <=  'sd153; // 726
        'h2d7: dout <=  'sd943; // 727
        'h2d8: dout <=  'sd2048; // 728
        'h2d9: dout <=  'sd1834; // 729
        'h2da: dout <= -'sd1407; // 730
        'h2db: dout <=  'sd1432; // 731
        'h2dc: dout <= -'sd1722; // 732
        'h2dd: dout <=  'sd897; // 733
        'h2de: dout <= -'sd978; // 734
        'h2df: dout <=  'sd2196; // 735
        'h2e0: dout <=  'sd953; // 736
        'h2e1: dout <= -'sd813; // 737
        'h2e2: dout <=  'sd1442; // 738
        'h2e3: dout <=  'sd2116; // 739
        'h2e4: dout <= -'sd424; // 740
        'h2e5: dout <= -'sd12; // 741
        'h2e6: dout <=  'sd945; // 742
        'h2e7: dout <= -'sd1149; // 743
        'h2e8: dout <= -'sd2181; // 744
        'h2e9: dout <= -'sd1370; // 745
        'h2ea: dout <=  'sd2063; // 746
        'h2eb: dout <=  'sd2138; // 747
        'h2ec: dout <=  'sd544; // 748
        'h2ed: dout <=  'sd666; // 749
        'h2ee: dout <=  'sd46; // 750
        'h2ef: dout <= -'sd1204; // 751
        'h2f0: dout <= -'sd1374; // 752
        'h2f1: dout <= -'sd672; // 753
        'h2f2: dout <=  'sd1177; // 754
        'h2f3: dout <=  'sd1601; // 755
        'h2f4: dout <=  'sd1255; // 756
        'h2f5: dout <=  'sd389; // 757
        'h2f6: dout <=  'sd1521; // 758
        'h2f7: dout <=  'sd767; // 759
        'h2f8: dout <= -'sd401; // 760
        'h2f9: dout <= -'sd1874; // 761
        'h2fa: dout <= -'sd1061; // 762
        'h2fb: dout <=  'sd2131; // 763
        'h2fc: dout <= -'sd654; // 764
        'h2fd: dout <= -'sd281; // 765
        'h2fe: dout <=  'sd621; // 766
        'h2ff: dout <= -'sd558; // 767
        'h300: dout <=  'sd22; // 768
        'h301: dout <= -'sd2209; // 769
        'h302: dout <= -'sd2218; // 770
        'h303: dout <=  'sd1173; // 771
        'h304: dout <= -'sd1761; // 772
        'h305: dout <=  'sd670; // 773
        'h306: dout <=  'sd1371; // 774
        'h307: dout <= -'sd485; // 775
        'h308: dout <= -'sd1928; // 776
        'h309: dout <= -'sd2014; // 777
        'h30a: dout <= -'sd2273; // 778
        'h30b: dout <= -'sd1003; // 779
        'h30c: dout <=  'sd1529; // 780
        'h30d: dout <= -'sd270; // 781
        'h30e: dout <= -'sd1879; // 782
        'h30f: dout <= -'sd1357; // 783
        'h310: dout <=  'sd1419; // 784
        'h311: dout <=  'sd2082; // 785
        'h312: dout <=  'sd386; // 786
        'h313: dout <=  'sd1947; // 787
        'h314: dout <=  'sd1553; // 788
        'h315: dout <= -'sd2036; // 789
        'h316: dout <=  'sd779; // 790
        'h317: dout <= -'sd651; // 791
        'h318: dout <=  'sd246; // 792
        'h319: dout <=  'sd863; // 793
        'h31a: dout <= -'sd942; // 794
        'h31b: dout <= -'sd803; // 795
        'h31c: dout <= -'sd645; // 796
        'h31d: dout <=  'sd486; // 797
        'h31e: dout <=  'sd1571; // 798
        'h31f: dout <= -'sd2099; // 799
        'h320: dout <= -'sd79; // 800
        'h321: dout <= -'sd1982; // 801
        'h322: dout <= -'sd2119; // 802
        'h323: dout <=  'sd1277; // 803
        'h324: dout <= -'sd1552; // 804
        'h325: dout <=  'sd1110; // 805
        'h326: dout <= -'sd2094; // 806
        'h327: dout <= -'sd1533; // 807
        'h328: dout <= -'sd981; // 808
        'h329: dout <=  'sd2006; // 809
        'h32a: dout <=  'sd1230; // 810
        'h32b: dout <= -'sd603; // 811
        'h32c: dout <=  'sd1509; // 812
        'h32d: dout <= -'sd1942; // 813
        'h32e: dout <=  'sd604; // 814
        'h32f: dout <=  'sd1620; // 815
        'h330: dout <=  'sd1405; // 816
        'h331: dout <= -'sd139; // 817
        'h332: dout <=  'sd726; // 818
        'h333: dout <= -'sd2060; // 819
        'h334: dout <=  'sd129; // 820
        'h335: dout <= -'sd1277; // 821
        'h336: dout <=  'sd183; // 822
        'h337: dout <= -'sd205; // 823
        'h338: dout <= -'sd1489; // 824
        'h339: dout <=  'sd2015; // 825
        'h33a: dout <= -'sd2225; // 826
        'h33b: dout <= -'sd1838; // 827
        'h33c: dout <=  'sd542; // 828
        'h33d: dout <=  'sd1854; // 829
        'h33e: dout <=  'sd1817; // 830
        'h33f: dout <=  'sd1531; // 831
        'h340: dout <=  'sd1550; // 832
        'h341: dout <= -'sd1708; // 833
        'h342: dout <= -'sd409; // 834
        'h343: dout <=  'sd63; // 835
        'h344: dout <= -'sd611; // 836
        'h345: dout <=  'sd408; // 837
        'h346: dout <= -'sd983; // 838
        'h347: dout <=  'sd709; // 839
        'h348: dout <= -'sd986; // 840
        'h349: dout <=  'sd1537; // 841
        'h34a: dout <= -'sd599; // 842
        'h34b: dout <= -'sd37; // 843
        'h34c: dout <=  'sd1588; // 844
        'h34d: dout <= -'sd155; // 845
        'h34e: dout <= -'sd898; // 846
        'h34f: dout <= -'sd2055; // 847
        'h350: dout <= -'sd1138; // 848
        'h351: dout <= -'sd1272; // 849
        'h352: dout <=  'sd22; // 850
        'h353: dout <=  'sd825; // 851
        'h354: dout <= -'sd493; // 852
        'h355: dout <= -'sd1968; // 853
        'h356: dout <= -'sd393; // 854
        'h357: dout <=  'sd1649; // 855
        'h358: dout <=  'sd420; // 856
        'h359: dout <=  'sd2254; // 857
        'h35a: dout <=  'sd1530; // 858
        'h35b: dout <=  'sd2151; // 859
        'h35c: dout <=  'sd1983; // 860
        'h35d: dout <=  'sd102; // 861
        'h35e: dout <= -'sd365; // 862
        'h35f: dout <= -'sd1925; // 863
        'h360: dout <=  'sd1033; // 864
        'h361: dout <=  'sd1773; // 865
        'h362: dout <=  'sd1465; // 866
        'h363: dout <=  'sd1934; // 867
        'h364: dout <=  'sd464; // 868
        'h365: dout <= -'sd1371; // 869
        'h366: dout <= -'sd1622; // 870
        'h367: dout <= -'sd1219; // 871
        'h368: dout <=  'sd810; // 872
        'h369: dout <= -'sd91; // 873
        'h36a: dout <= -'sd1110; // 874
        'h36b: dout <= -'sd256; // 875
        'h36c: dout <= -'sd1091; // 876
        'h36d: dout <= -'sd148; // 877
        'h36e: dout <=  'sd1792; // 878
        'h36f: dout <=  'sd823; // 879
        'h370: dout <=  'sd1431; // 880
        'h371: dout <= -'sd412; // 881
        'h372: dout <= -'sd135; // 882
        'h373: dout <= -'sd1871; // 883
        'h374: dout <= -'sd255; // 884
        'h375: dout <=  'sd2165; // 885
        'h376: dout <= -'sd362; // 886
        'h377: dout <= -'sd56; // 887
        'h378: dout <=  'sd1610; // 888
        'h379: dout <=  'sd2162; // 889
        'h37a: dout <= -'sd938; // 890
        'h37b: dout <=  'sd1537; // 891
        'h37c: dout <=  'sd180; // 892
        'h37d: dout <= -'sd841; // 893
        'h37e: dout <= -'sd1680; // 894
        'h37f: dout <= -'sd139; // 895
        'h380: dout <= -'sd1121; // 896
        'h381: dout <=  'sd2291; // 897
        'h382: dout <= -'sd969; // 898
        'h383: dout <= -'sd1752; // 899
        'h384: dout <= -'sd467; // 900
        'h385: dout <=  'sd281; // 901
        'h386: dout <= -'sd2096; // 902
        'h387: dout <=  'sd330; // 903
        'h388: dout <= -'sd2275; // 904
        'h389: dout <=  'sd1185; // 905
        'h38a: dout <= -'sd662; // 906
        'h38b: dout <=  'sd1545; // 907
        'h38c: dout <= -'sd447; // 908
        'h38d: dout <=  'sd2114; // 909
        'h38e: dout <=  'sd164; // 910
        'h38f: dout <=  'sd716; // 911
        'h390: dout <= -'sd786; // 912
        'h391: dout <=  'sd2003; // 913
        'h392: dout <=  'sd379; // 914
        'h393: dout <=  'sd970; // 915
        'h394: dout <=  'sd445; // 916
        'h395: dout <= -'sd290; // 917
        'h396: dout <= -'sd2160; // 918
        'h397: dout <=  'sd1668; // 919
        'h398: dout <=  'sd1410; // 920
        'h399: dout <=  'sd1371; // 921
        'h39a: dout <= -'sd1413; // 922
        'h39b: dout <=  'sd1416; // 923
        'h39c: dout <=  'sd807; // 924
        'h39d: dout <=  'sd771; // 925
        'h39e: dout <= -'sd692; // 926
        'h39f: dout <=  'sd1587; // 927
        'h3a0: dout <= -'sd1514; // 928
        'h3a1: dout <=  'sd561; // 929
        'h3a2: dout <= -'sd2210; // 930
        'h3a3: dout <= -'sd788; // 931
        'h3a4: dout <= -'sd243; // 932
        'h3a5: dout <=  'sd443; // 933
        'h3a6: dout <=  'sd305; // 934
        'h3a7: dout <=  'sd256; // 935
        'h3a8: dout <=  'sd1701; // 936
        'h3a9: dout <= -'sd1532; // 937
        'h3aa: dout <=  'sd113; // 938
        'h3ab: dout <=  'sd1563; // 939
        'h3ac: dout <= -'sd1490; // 940
        'h3ad: dout <= -'sd319; // 941
        'h3ae: dout <=  'sd1640; // 942
        'h3af: dout <=  'sd2160; // 943
        'h3b0: dout <= -'sd498; // 944
        'h3b1: dout <=  'sd677; // 945
        'h3b2: dout <=  'sd1097; // 946
        'h3b3: dout <= -'sd1081; // 947
        'h3b4: dout <= -'sd1251; // 948
        'h3b5: dout <=  'sd1429; // 949
        'h3b6: dout <=  'sd2024; // 950
        'h3b7: dout <= -'sd9; // 951
        'h3b8: dout <=  'sd1107; // 952
        'h3b9: dout <= -'sd1591; // 953
        'h3ba: dout <=  'sd849; // 954
        'h3bb: dout <= -'sd191; // 955
        'h3bc: dout <=  'sd1325; // 956
        'h3bd: dout <= -'sd1256; // 957
        'h3be: dout <=  'sd110; // 958
        'h3bf: dout <=  'sd918; // 959
        'h3c0: dout <=  'sd1694; // 960
        'h3c1: dout <= -'sd1103; // 961
        'h3c2: dout <= -'sd750; // 962
        'h3c3: dout <= -'sd124; // 963
        'h3c4: dout <=  'sd491; // 964
        'h3c5: dout <=  'sd762; // 965
        'h3c6: dout <= -'sd2206; // 966
        'h3c7: dout <= -'sd1287; // 967
        'h3c8: dout <=  'sd584; // 968
        'h3c9: dout <= -'sd1301; // 969
        'h3ca: dout <=  'sd477; // 970
        'h3cb: dout <= -'sd1868; // 971
        'h3cc: dout <=  'sd2187; // 972
        'h3cd: dout <=  'sd76; // 973
        'h3ce: dout <=  'sd2110; // 974
        'h3cf: dout <=  'sd1633; // 975
        'h3d0: dout <=  'sd274; // 976
        'h3d1: dout <= -'sd885; // 977
        'h3d2: dout <=  'sd2246; // 978
        'h3d3: dout <= -'sd606; // 979
        'h3d4: dout <=  'sd645; // 980
        'h3d5: dout <= -'sd1378; // 981
        'h3d6: dout <=  'sd237; // 982
        'h3d7: dout <=  'sd433; // 983
        'h3d8: dout <=  'sd1255; // 984
        'h3d9: dout <= -'sd82; // 985
        'h3da: dout <=  'sd1129; // 986
        'h3db: dout <= -'sd34; // 987
        'h3dc: dout <=  'sd144; // 988
        'h3dd: dout <=  'sd80; // 989
        'h3de: dout <= -'sd827; // 990
        'h3df: dout <=  'sd803; // 991
        'h3e0: dout <=  'sd1809; // 992
        'h3e1: dout <= -'sd1369; // 993
        'h3e2: dout <=  'sd250; // 994
        'h3e3: dout <=  'sd184; // 995
        'h3e4: dout <=  'sd1368; // 996
        'h3e5: dout <= -'sd486; // 997
        'h3e6: dout <= -'sd2069; // 998
        'h3e7: dout <=  'sd2126; // 999
        'h3e8: dout <= -'sd318; // 1000
        'h3e9: dout <=  'sd1946; // 1001
        'h3ea: dout <=  'sd2107; // 1002
        'h3eb: dout <= -'sd1969; // 1003
        'h3ec: dout <= -'sd64; // 1004
        'h3ed: dout <=  'sd2117; // 1005
        'h3ee: dout <= -'sd1762; // 1006
        'h3ef: dout <= -'sd945; // 1007
        'h3f0: dout <= -'sd1181; // 1008
        'h3f1: dout <=  'sd731; // 1009
        'h3f2: dout <= -'sd360; // 1010
        'h3f3: dout <= -'sd1804; // 1011
        'h3f4: dout <=  'sd1675; // 1012
        'h3f5: dout <=  'sd693; // 1013
        'h3f6: dout <=  'sd319; // 1014
        'h3f7: dout <=  'sd1638; // 1015
        'h3f8: dout <=  'sd1132; // 1016
        'h3f9: dout <=  'sd198; // 1017
        'h3fa: dout <=  'sd185; // 1018
        'h3fb: dout <=  'sd2236; // 1019
        'h3fc: dout <= -'sd1951; // 1020
        'h3fd: dout <= -'sd865; // 1021
        'h3fe: dout <= -'sd1098; // 1022
        'h3ff: dout <=  'sd145; // 1023
        'h400: dout <=  'sd816; // 1024
        'h401: dout <=  'sd353; // 1025
        'h402: dout <=  'sd1032; // 1026
        'h403: dout <= -'sd2114; // 1027
        'h404: dout <= -'sd1740; // 1028
        'h405: dout <= -'sd659; // 1029
        'h406: dout <= -'sd735; // 1030
        'h407: dout <=  'sd1307; // 1031
        'h408: dout <= -'sd156; // 1032
        'h409: dout <=  'sd1194; // 1033
        'h40a: dout <= -'sd1190; // 1034
        'h40b: dout <=  'sd215; // 1035
        'h40c: dout <= -'sd1918; // 1036
        'h40d: dout <=  'sd25; // 1037
        'h40e: dout <=  'sd1259; // 1038
        'h40f: dout <=  'sd1320; // 1039
        'h410: dout <= -'sd1074; // 1040
        'h411: dout <=  'sd1327; // 1041
        'h412: dout <=  'sd832; // 1042
        'h413: dout <= -'sd975; // 1043
        'h414: dout <= -'sd1299; // 1044
        'h415: dout <=  'sd392; // 1045
        'h416: dout <=  'sd321; // 1046
        'h417: dout <= -'sd576; // 1047
        'h418: dout <=  'sd152; // 1048
        'h419: dout <=  'sd1488; // 1049
        'h41a: dout <= -'sd1331; // 1050
        'h41b: dout <=  'sd938; // 1051
        'h41c: dout <= -'sd1174; // 1052
        'h41d: dout <= -'sd1399; // 1053
        'h41e: dout <= -'sd1487; // 1054
        'h41f: dout <= -'sd1113; // 1055
        'h420: dout <=  'sd1078; // 1056
        'h421: dout <=  'sd401; // 1057
        'h422: dout <=  'sd706; // 1058
        'h423: dout <= -'sd1792; // 1059
        'h424: dout <=  'sd1157; // 1060
        'h425: dout <=  'sd465; // 1061
        'h426: dout <= -'sd815; // 1062
        'h427: dout <= -'sd199; // 1063
        'h428: dout <=  'sd510; // 1064
        'h429: dout <=  'sd299; // 1065
        'h42a: dout <= -'sd2207; // 1066
        'h42b: dout <= -'sd686; // 1067
        'h42c: dout <=  'sd2128; // 1068
        'h42d: dout <=  'sd193; // 1069
        'h42e: dout <=  'sd1500; // 1070
        'h42f: dout <=  'sd2169; // 1071
        'h430: dout <= -'sd443; // 1072
        'h431: dout <= -'sd191; // 1073
        'h432: dout <=  'sd670; // 1074
        'h433: dout <= -'sd1880; // 1075
        'h434: dout <=  'sd2233; // 1076
        'h435: dout <= -'sd2056; // 1077
        'h436: dout <= -'sd1907; // 1078
        'h437: dout <= -'sd1337; // 1079
        'h438: dout <=  'sd825; // 1080
        'h439: dout <= -'sd213; // 1081
        'h43a: dout <=  'sd833; // 1082
        'h43b: dout <= -'sd1278; // 1083
        'h43c: dout <= -'sd369; // 1084
        'h43d: dout <= -'sd1499; // 1085
        'h43e: dout <=  'sd1650; // 1086
        'h43f: dout <= -'sd2044; // 1087
        'h440: dout <= -'sd57; // 1088
        'h441: dout <=  'sd334; // 1089
        'h442: dout <=  'sd162; // 1090
        'h443: dout <= -'sd2174; // 1091
        'h444: dout <= -'sd2044; // 1092
        'h445: dout <=  'sd1116; // 1093
        'h446: dout <= -'sd1838; // 1094
        'h447: dout <=  'sd990; // 1095
        'h448: dout <=  'sd1671; // 1096
        'h449: dout <=  'sd1082; // 1097
        'h44a: dout <= -'sd1680; // 1098
        'h44b: dout <=  'sd1089; // 1099
        'h44c: dout <=  'sd73; // 1100
        'h44d: dout <= -'sd293; // 1101
        'h44e: dout <=  'sd397; // 1102
        'h44f: dout <=  'sd426; // 1103
        'h450: dout <= -'sd104; // 1104
        'h451: dout <= -'sd1191; // 1105
        'h452: dout <=  'sd130; // 1106
        'h453: dout <= -'sd211; // 1107
        'h454: dout <= -'sd790; // 1108
        'h455: dout <= -'sd1070; // 1109
        'h456: dout <=  'sd1675; // 1110
        'h457: dout <= -'sd275; // 1111
        'h458: dout <= -'sd2130; // 1112
        'h459: dout <= -'sd1077; // 1113
        'h45a: dout <= -'sd870; // 1114
        'h45b: dout <= -'sd1081; // 1115
        'h45c: dout <= -'sd375; // 1116
        'h45d: dout <= -'sd1914; // 1117
        'h45e: dout <= -'sd1237; // 1118
        'h45f: dout <= -'sd1252; // 1119
        'h460: dout <= -'sd514; // 1120
        'h461: dout <=  'sd471; // 1121
        'h462: dout <=  'sd2142; // 1122
        'h463: dout <= -'sd1193; // 1123
        'h464: dout <=  'sd164; // 1124
        'h465: dout <=  'sd2043; // 1125
        'h466: dout <= -'sd2289; // 1126
        'h467: dout <=  'sd747; // 1127
        'h468: dout <=  'sd1629; // 1128
        'h469: dout <= -'sd636; // 1129
        'h46a: dout <=  'sd683; // 1130
        'h46b: dout <=  'sd134; // 1131
        'h46c: dout <= -'sd171; // 1132
        'h46d: dout <= -'sd802; // 1133
        'h46e: dout <=  'sd58; // 1134
        'h46f: dout <=  'sd2117; // 1135
        'h470: dout <=  'sd1173; // 1136
        'h471: dout <= -'sd1026; // 1137
        'h472: dout <=  'sd1931; // 1138
        'h473: dout <=  'sd2159; // 1139
        'h474: dout <=  'sd1710; // 1140
        'h475: dout <=  'sd485; // 1141
        'h476: dout <=  'sd989; // 1142
        'h477: dout <=  'sd1479; // 1143
        'h478: dout <=  'sd649; // 1144
        'h479: dout <= -'sd1921; // 1145
        'h47a: dout <=  'sd1488; // 1146
        'h47b: dout <=  'sd790; // 1147
        'h47c: dout <=  'sd53; // 1148
        'h47d: dout <=  'sd1997; // 1149
        'h47e: dout <= -'sd1687; // 1150
        'h47f: dout <=  'sd2063; // 1151
        'h480: dout <=  'sd1803; // 1152
        'h481: dout <= -'sd2; // 1153
        'h482: dout <= -'sd745; // 1154
        'h483: dout <=  'sd1472; // 1155
        'h484: dout <= -'sd914; // 1156
        'h485: dout <=  'sd790; // 1157
        'h486: dout <= -'sd1064; // 1158
        'h487: dout <=  'sd116; // 1159
        'h488: dout <= -'sd2249; // 1160
        'h489: dout <= -'sd589; // 1161
        'h48a: dout <= -'sd541; // 1162
        'h48b: dout <= -'sd1100; // 1163
        'h48c: dout <=  'sd1079; // 1164
        'h48d: dout <=  'sd1236; // 1165
        'h48e: dout <=  'sd1118; // 1166
        'h48f: dout <=  'sd1523; // 1167
        'h490: dout <= -'sd1187; // 1168
        'h491: dout <=  'sd1242; // 1169
        'h492: dout <= -'sd1548; // 1170
        'h493: dout <= -'sd1769; // 1171
        'h494: dout <= -'sd40; // 1172
        'h495: dout <= -'sd1772; // 1173
        'h496: dout <=  'sd1657; // 1174
        'h497: dout <=  'sd279; // 1175
        'h498: dout <=  'sd1081; // 1176
        'h499: dout <=  'sd1653; // 1177
        'h49a: dout <=  'sd1815; // 1178
        'h49b: dout <=  'sd1553; // 1179
        'h49c: dout <= -'sd639; // 1180
        'h49d: dout <=  'sd1158; // 1181
        'h49e: dout <=  'sd14; // 1182
        'h49f: dout <= -'sd711; // 1183
        'h4a0: dout <=  'sd936; // 1184
        'h4a1: dout <= -'sd1043; // 1185
        'h4a2: dout <= -'sd65; // 1186
        'h4a3: dout <=  'sd1843; // 1187
        'h4a4: dout <=  'sd1876; // 1188
        'h4a5: dout <= -'sd807; // 1189
        'h4a6: dout <=  'sd1102; // 1190
        'h4a7: dout <=  'sd926; // 1191
        'h4a8: dout <= -'sd839; // 1192
        'h4a9: dout <= -'sd1603; // 1193
        'h4aa: dout <=  'sd179; // 1194
        'h4ab: dout <=  'sd1630; // 1195
        'h4ac: dout <=  'sd2152; // 1196
        'h4ad: dout <= -'sd1021; // 1197
        'h4ae: dout <=  'sd908; // 1198
        'h4af: dout <= -'sd1435; // 1199
        'h4b0: dout <=  'sd2251; // 1200
        'h4b1: dout <=  'sd76; // 1201
        'h4b2: dout <= -'sd572; // 1202
        'h4b3: dout <= -'sd1151; // 1203
        'h4b4: dout <=  'sd1735; // 1204
        'h4b5: dout <=  'sd686; // 1205
        'h4b6: dout <=  'sd897; // 1206
        'h4b7: dout <=  'sd2227; // 1207
        'h4b8: dout <= -'sd1518; // 1208
        'h4b9: dout <=  'sd2171; // 1209
        'h4ba: dout <=  'sd1065; // 1210
        'h4bb: dout <=  'sd307; // 1211
        'h4bc: dout <= -'sd1810; // 1212
        'h4bd: dout <=  'sd664; // 1213
        'h4be: dout <=  'sd2248; // 1214
        'h4bf: dout <=  'sd1618; // 1215
        'h4c0: dout <= -'sd689; // 1216
        'h4c1: dout <= -'sd1856; // 1217
        'h4c2: dout <= -'sd148; // 1218
        'h4c3: dout <= -'sd758; // 1219
        'h4c4: dout <= -'sd1989; // 1220
        'h4c5: dout <= -'sd242; // 1221
        'h4c6: dout <= -'sd1528; // 1222
        'h4c7: dout <=  'sd1304; // 1223
        'h4c8: dout <=  'sd1115; // 1224
        'h4c9: dout <=  'sd258; // 1225
        'h4ca: dout <= -'sd1457; // 1226
        'h4cb: dout <=  'sd2213; // 1227
        'h4cc: dout <=  'sd1936; // 1228
        'h4cd: dout <= -'sd1577; // 1229
        'h4ce: dout <= -'sd1504; // 1230
        'h4cf: dout <= -'sd1502; // 1231
        'h4d0: dout <=  'sd698; // 1232
        'h4d1: dout <=  'sd2055; // 1233
        'h4d2: dout <=  'sd536; // 1234
        'h4d3: dout <=  'sd1988; // 1235
        'h4d4: dout <= -'sd2153; // 1236
        'h4d5: dout <=  'sd1737; // 1237
        'h4d6: dout <=  'sd2134; // 1238
        'h4d7: dout <= -'sd1005; // 1239
        'h4d8: dout <= -'sd294; // 1240
        'h4d9: dout <= -'sd404; // 1241
        'h4da: dout <= -'sd2049; // 1242
        'h4db: dout <= -'sd329; // 1243
        'h4dc: dout <= -'sd473; // 1244
        'h4dd: dout <=  'sd1626; // 1245
        'h4de: dout <= -'sd685; // 1246
        'h4df: dout <=  'sd73; // 1247
        'h4e0: dout <=  'sd926; // 1248
        'h4e1: dout <= -'sd2247; // 1249
        'h4e2: dout <=  'sd309; // 1250
        'h4e3: dout <=  'sd932; // 1251
        'h4e4: dout <=  'sd1524; // 1252
        'h4e5: dout <=  'sd1944; // 1253
        'h4e6: dout <=  'sd1446; // 1254
        'h4e7: dout <= -'sd123; // 1255
        'h4e8: dout <= -'sd502; // 1256
        'h4e9: dout <= -'sd1519; // 1257
        'h4ea: dout <=  'sd1980; // 1258
        'h4eb: dout <=  'sd1270; // 1259
        'h4ec: dout <= -'sd1835; // 1260
        'h4ed: dout <= -'sd1977; // 1261
        'h4ee: dout <=  'sd2194; // 1262
        'h4ef: dout <= -'sd1826; // 1263
        'h4f0: dout <= -'sd2046; // 1264
        'h4f1: dout <= -'sd2253; // 1265
        'h4f2: dout <=  'sd1641; // 1266
        'h4f3: dout <=  'sd1007; // 1267
        'h4f4: dout <=  'sd524; // 1268
        'h4f5: dout <=  'sd186; // 1269
        'h4f6: dout <= -'sd7; // 1270
        'h4f7: dout <=  'sd768; // 1271
        'h4f8: dout <=  'sd1962; // 1272
        'h4f9: dout <= -'sd1538; // 1273
        'h4fa: dout <=  'sd630; // 1274
        'h4fb: dout <= -'sd1466; // 1275
        'h4fc: dout <=  'sd272; // 1276
        'h4fd: dout <= -'sd1762; // 1277
        'h4fe: dout <= -'sd343; // 1278
        'h4ff: dout <=  'sd1012; // 1279
        'h500: dout <= -'sd1872; // 1280
        'h501: dout <=  'sd752; // 1281
        'h502: dout <= -'sd2004; // 1282
        'h503: dout <= -'sd1854; // 1283
        'h504: dout <= -'sd441; // 1284
        'h505: dout <=  'sd2249; // 1285
        'h506: dout <=  'sd912; // 1286
        'h507: dout <= -'sd1344; // 1287
        'h508: dout <=  'sd315; // 1288
        'h509: dout <= -'sd1437; // 1289
        'h50a: dout <= -'sd1099; // 1290
        'h50b: dout <= -'sd1359; // 1291
        'h50c: dout <= -'sd864; // 1292
        'h50d: dout <=  'sd272; // 1293
        'h50e: dout <=  'sd1483; // 1294
        'h50f: dout <=  'sd761; // 1295
        'h510: dout <=  'sd1539; // 1296
        'h511: dout <=  'sd63; // 1297
        'h512: dout <=  'sd852; // 1298
        'h513: dout <=  'sd1125; // 1299
        'h514: dout <=  'sd204; // 1300
        'h515: dout <= -'sd1376; // 1301
        'h516: dout <= -'sd1115; // 1302
        'h517: dout <= -'sd1794; // 1303
        'h518: dout <=  'sd1907; // 1304
        'h519: dout <= -'sd144; // 1305
        'h51a: dout <= -'sd132; // 1306
        'h51b: dout <=  'sd1751; // 1307
        'h51c: dout <=  'sd613; // 1308
        'h51d: dout <=  'sd10; // 1309
        'h51e: dout <= -'sd364; // 1310
        'h51f: dout <= -'sd2288; // 1311
        'h520: dout <=  'sd1362; // 1312
        'h521: dout <= -'sd144; // 1313
        'h522: dout <= -'sd1772; // 1314
        'h523: dout <=  'sd986; // 1315
        'h524: dout <= -'sd1485; // 1316
        'h525: dout <= -'sd298; // 1317
        'h526: dout <= -'sd143; // 1318
        'h527: dout <=  'sd2039; // 1319
        'h528: dout <=  'sd643; // 1320
        'h529: dout <= -'sd538; // 1321
        'h52a: dout <= -'sd1463; // 1322
        'h52b: dout <=  'sd359; // 1323
        'h52c: dout <= -'sd1679; // 1324
        'h52d: dout <=  'sd614; // 1325
        'h52e: dout <=  'sd1327; // 1326
        'h52f: dout <=  'sd998; // 1327
        'h530: dout <=  'sd771; // 1328
        'h531: dout <=  'sd788; // 1329
        'h532: dout <=  'sd1605; // 1330
        'h533: dout <= -'sd745; // 1331
        'h534: dout <= -'sd1665; // 1332
        'h535: dout <= -'sd1159; // 1333
        'h536: dout <= -'sd2025; // 1334
        'h537: dout <=  'sd1173; // 1335
        'h538: dout <=  'sd1118; // 1336
        'h539: dout <= -'sd427; // 1337
        'h53a: dout <= -'sd118; // 1338
        'h53b: dout <= -'sd1223; // 1339
        'h53c: dout <= -'sd1751; // 1340
        'h53d: dout <=  'sd1783; // 1341
        'h53e: dout <= -'sd332; // 1342
        'h53f: dout <= -'sd2127; // 1343
        'h540: dout <=  'sd574; // 1344
        'h541: dout <= -'sd1980; // 1345
        'h542: dout <=  'sd1440; // 1346
        'h543: dout <=  'sd949; // 1347
        'h544: dout <=  'sd2019; // 1348
        'h545: dout <=  'sd2005; // 1349
        'h546: dout <= -'sd805; // 1350
        'h547: dout <=  'sd594; // 1351
        'h548: dout <= -'sd2289; // 1352
        'h549: dout <= -'sd941; // 1353
        'h54a: dout <= -'sd1017; // 1354
        'h54b: dout <=  'sd1672; // 1355
        'h54c: dout <= -'sd266; // 1356
        'h54d: dout <=  'sd421; // 1357
        'h54e: dout <= -'sd1065; // 1358
        'h54f: dout <= -'sd169; // 1359
        'h550: dout <=  'sd1191; // 1360
        'h551: dout <= -'sd922; // 1361
        'h552: dout <=  'sd1922; // 1362
        'h553: dout <= -'sd1997; // 1363
        'h554: dout <=  'sd355; // 1364
        'h555: dout <= -'sd790; // 1365
        'h556: dout <=  'sd2097; // 1366
        'h557: dout <=  'sd1128; // 1367
        'h558: dout <=  'sd1376; // 1368
        'h559: dout <=  'sd1765; // 1369
        'h55a: dout <=  'sd1938; // 1370
        'h55b: dout <=  'sd595; // 1371
        'h55c: dout <=  'sd1734; // 1372
        'h55d: dout <=  'sd2156; // 1373
        'h55e: dout <=  'sd2162; // 1374
        'h55f: dout <=  'sd1962; // 1375
        'h560: dout <= -'sd1216; // 1376
        'h561: dout <=  'sd851; // 1377
        'h562: dout <= -'sd675; // 1378
        'h563: dout <= -'sd642; // 1379
        'h564: dout <=  'sd1140; // 1380
        'h565: dout <= -'sd187; // 1381
        'h566: dout <= -'sd1552; // 1382
        'h567: dout <= -'sd1965; // 1383
        'h568: dout <=  'sd1178; // 1384
        'h569: dout <=  'sd633; // 1385
        'h56a: dout <= -'sd1094; // 1386
        'h56b: dout <= -'sd2064; // 1387
        'h56c: dout <= -'sd2006; // 1388
        'h56d: dout <= -'sd1834; // 1389
        'h56e: dout <= -'sd1524; // 1390
        'h56f: dout <=  'sd2051; // 1391
        'h570: dout <=  'sd1690; // 1392
        'h571: dout <= -'sd2198; // 1393
        'h572: dout <= -'sd1231; // 1394
        'h573: dout <= -'sd2205; // 1395
        'h574: dout <=  'sd586; // 1396
        'h575: dout <= -'sd1244; // 1397
        'h576: dout <=  'sd1718; // 1398
        'h577: dout <=  'sd1232; // 1399
        'h578: dout <= -'sd724; // 1400
        'h579: dout <= -'sd1766; // 1401
        'h57a: dout <=  'sd1086; // 1402
        'h57b: dout <= -'sd478; // 1403
        'h57c: dout <= -'sd930; // 1404
        'h57d: dout <= -'sd2193; // 1405
        'h57e: dout <= -'sd2238; // 1406
        'h57f: dout <=  'sd250; // 1407
        'h580: dout <= -'sd2253; // 1408
        'h581: dout <= -'sd1415; // 1409
        'h582: dout <= -'sd722; // 1410
        'h583: dout <=  'sd1868; // 1411
        'h584: dout <=  'sd1930; // 1412
        'h585: dout <=  'sd1917; // 1413
        'h586: dout <= -'sd1098; // 1414
        'h587: dout <=  'sd612; // 1415
        'h588: dout <=  'sd88; // 1416
        'h589: dout <= -'sd228; // 1417
        'h58a: dout <= -'sd28; // 1418
        'h58b: dout <=  'sd2153; // 1419
        'h58c: dout <=  'sd1424; // 1420
        'h58d: dout <=  'sd105; // 1421
        'h58e: dout <=  'sd1840; // 1422
        'h58f: dout <= -'sd2211; // 1423
        'h590: dout <=  'sd1079; // 1424
        'h591: dout <=  'sd823; // 1425
        'h592: dout <= -'sd1008; // 1426
        'h593: dout <= -'sd340; // 1427
        'h594: dout <= -'sd1725; // 1428
        'h595: dout <= -'sd1874; // 1429
        'h596: dout <= -'sd919; // 1430
        'h597: dout <= -'sd598; // 1431
        'h598: dout <= -'sd467; // 1432
        'h599: dout <= -'sd2107; // 1433
        'h59a: dout <=  'sd1862; // 1434
        'h59b: dout <= -'sd860; // 1435
        'h59c: dout <=  'sd154; // 1436
        'h59d: dout <= -'sd557; // 1437
        'h59e: dout <= -'sd235; // 1438
        'h59f: dout <=  'sd2169; // 1439
        'h5a0: dout <= -'sd1089; // 1440
        'h5a1: dout <= -'sd107; // 1441
        'h5a2: dout <=  'sd1210; // 1442
        'h5a3: dout <= -'sd1139; // 1443
        'h5a4: dout <=  'sd1663; // 1444
        'h5a5: dout <= -'sd673; // 1445
        'h5a6: dout <= -'sd1959; // 1446
        'h5a7: dout <=  'sd1943; // 1447
        'h5a8: dout <= -'sd963; // 1448
        'h5a9: dout <=  'sd984; // 1449
        'h5aa: dout <=  'sd2091; // 1450
        'h5ab: dout <=  'sd2020; // 1451
        'h5ac: dout <=  'sd1238; // 1452
        'h5ad: dout <= -'sd1; // 1453
        'h5ae: dout <= -'sd520; // 1454
        'h5af: dout <= -'sd897; // 1455
        'h5b0: dout <= -'sd609; // 1456
        'h5b1: dout <= -'sd165; // 1457
        'h5b2: dout <=  'sd1669; // 1458
        'h5b3: dout <= -'sd1768; // 1459
        'h5b4: dout <= -'sd2186; // 1460
        'h5b5: dout <=  'sd1367; // 1461
        'h5b6: dout <=  'sd623; // 1462
        'h5b7: dout <=  'sd2118; // 1463
        'h5b8: dout <= -'sd681; // 1464
        'h5b9: dout <= -'sd1912; // 1465
        'h5ba: dout <=  'sd254; // 1466
        'h5bb: dout <= -'sd1167; // 1467
        'h5bc: dout <= -'sd2090; // 1468
        'h5bd: dout <=  'sd861; // 1469
        'h5be: dout <= -'sd1301; // 1470
        'h5bf: dout <= -'sd327; // 1471
        'h5c0: dout <=  'sd1859; // 1472
        'h5c1: dout <=  'sd28; // 1473
        'h5c2: dout <= -'sd34; // 1474
        'h5c3: dout <=  'sd2219; // 1475
        'h5c4: dout <= -'sd1161; // 1476
        'h5c5: dout <= -'sd2097; // 1477
        'h5c6: dout <=  'sd2045; // 1478
        'h5c7: dout <= -'sd1133; // 1479
        'h5c8: dout <= -'sd697; // 1480
        'h5c9: dout <= -'sd2194; // 1481
        'h5ca: dout <= -'sd735; // 1482
        'h5cb: dout <=  'sd853; // 1483
        'h5cc: dout <= -'sd345; // 1484
        'h5cd: dout <=  'sd660; // 1485
        'h5ce: dout <=  'sd984; // 1486
        'h5cf: dout <=  'sd2216; // 1487
        'h5d0: dout <= -'sd2229; // 1488
        'h5d1: dout <= -'sd317; // 1489
        'h5d2: dout <= -'sd71; // 1490
        'h5d3: dout <=  'sd234; // 1491
        'h5d4: dout <= -'sd1915; // 1492
        'h5d5: dout <=  'sd2070; // 1493
        'h5d6: dout <= -'sd1380; // 1494
        'h5d7: dout <= -'sd1902; // 1495
        'h5d8: dout <=  'sd1617; // 1496
        'h5d9: dout <= -'sd217; // 1497
        'h5da: dout <= -'sd663; // 1498
        'h5db: dout <= -'sd398; // 1499
        'h5dc: dout <= -'sd737; // 1500
        'h5dd: dout <=  'sd2275; // 1501
        'h5de: dout <= -'sd1458; // 1502
        'h5df: dout <=  'sd415; // 1503
        'h5e0: dout <=  'sd1515; // 1504
        'h5e1: dout <=  'sd427; // 1505
        'h5e2: dout <= -'sd1739; // 1506
        'h5e3: dout <=  'sd1903; // 1507
        'h5e4: dout <=  'sd619; // 1508
        'h5e5: dout <=  'sd2193; // 1509
        'h5e6: dout <=  'sd446; // 1510
        'h5e7: dout <= -'sd473; // 1511
        'h5e8: dout <=  'sd1209; // 1512
        'h5e9: dout <=  'sd805; // 1513
        'h5ea: dout <= -'sd1838; // 1514
        'h5eb: dout <=  'sd1009; // 1515
        'h5ec: dout <= -'sd820; // 1516
        'h5ed: dout <= -'sd1850; // 1517
        'h5ee: dout <= -'sd986; // 1518
        'h5ef: dout <=  'sd1355; // 1519
        'h5f0: dout <=  'sd992; // 1520
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hp_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <= -'sd456; // 0
        'h001: dout <= -'sd912; // 1
        'h002: dout <=  'sd1248; // 2
        'h003: dout <= -'sd133; // 3
        'h004: dout <= -'sd441; // 4
        'h005: dout <= -'sd1508; // 5
        'h006: dout <=  'sd2102; // 6
        'h007: dout <= -'sd194; // 7
        'h008: dout <= -'sd22; // 8
        'h009: dout <= -'sd226; // 9
        'h00a: dout <=  'sd732; // 10
        'h00b: dout <=  'sd1480; // 11
        'h00c: dout <=  'sd596; // 12
        'h00d: dout <= -'sd396; // 13
        'h00e: dout <= -'sd2202; // 14
        'h00f: dout <= -'sd1337; // 15
        'h010: dout <= -'sd823; // 16
        'h011: dout <=  'sd1239; // 17
        'h012: dout <=  'sd1932; // 18
        'h013: dout <= -'sd936; // 19
        'h014: dout <= -'sd1161; // 20
        'h015: dout <=  'sd722; // 21
        'h016: dout <=  'sd101; // 22
        'h017: dout <=  'sd2069; // 23
        'h018: dout <= -'sd273; // 24
        'h019: dout <= -'sd2155; // 25
        'h01a: dout <=  'sd1729; // 26
        'h01b: dout <=  'sd1042; // 27
        'h01c: dout <= -'sd1849; // 28
        'h01d: dout <=  'sd2236; // 29
        'h01e: dout <= -'sd254; // 30
        'h01f: dout <=  'sd2114; // 31
        'h020: dout <=  'sd1525; // 32
        'h021: dout <=  'sd138; // 33
        'h022: dout <=  'sd1693; // 34
        'h023: dout <= -'sd1800; // 35
        'h024: dout <= -'sd1420; // 36
        'h025: dout <=  'sd471; // 37
        'h026: dout <= -'sd273; // 38
        'h027: dout <=  'sd1723; // 39
        'h028: dout <= -'sd278; // 40
        'h029: dout <=  'sd172; // 41
        'h02a: dout <=  'sd2008; // 42
        'h02b: dout <= -'sd1181; // 43
        'h02c: dout <= -'sd427; // 44
        'h02d: dout <=  'sd1566; // 45
        'h02e: dout <= -'sd1891; // 46
        'h02f: dout <=  'sd681; // 47
        'h030: dout <= -'sd408; // 48
        'h031: dout <= -'sd865; // 49
        'h032: dout <=  'sd5; // 50
        'h033: dout <= -'sd1022; // 51
        'h034: dout <= -'sd1073; // 52
        'h035: dout <=  'sd2223; // 53
        'h036: dout <= -'sd1645; // 54
        'h037: dout <=  'sd2165; // 55
        'h038: dout <= -'sd1952; // 56
        'h039: dout <=  'sd1690; // 57
        'h03a: dout <= -'sd1916; // 58
        'h03b: dout <=  'sd1742; // 59
        'h03c: dout <= -'sd346; // 60
        'h03d: dout <=  'sd668; // 61
        'h03e: dout <=  'sd1062; // 62
        'h03f: dout <= -'sd42; // 63
        'h040: dout <=  'sd774; // 64
        'h041: dout <=  'sd67; // 65
        'h042: dout <=  'sd1472; // 66
        'h043: dout <= -'sd1836; // 67
        'h044: dout <= -'sd2276; // 68
        'h045: dout <=  'sd1882; // 69
        'h046: dout <= -'sd1930; // 70
        'h047: dout <=  'sd542; // 71
        'h048: dout <= -'sd756; // 72
        'h049: dout <= -'sd697; // 73
        'h04a: dout <=  'sd1618; // 74
        'h04b: dout <= -'sd159; // 75
        'h04c: dout <= -'sd561; // 76
        'h04d: dout <=  'sd936; // 77
        'h04e: dout <= -'sd1143; // 78
        'h04f: dout <=  'sd1277; // 79
        'h050: dout <= -'sd292; // 80
        'h051: dout <=  'sd874; // 81
        'h052: dout <= -'sd411; // 82
        'h053: dout <=  'sd263; // 83
        'h054: dout <=  'sd133; // 84
        'h055: dout <=  'sd1475; // 85
        'h056: dout <=  'sd403; // 86
        'h057: dout <= -'sd1510; // 87
        'h058: dout <=  'sd431; // 88
        'h059: dout <= -'sd1216; // 89
        'h05a: dout <=  'sd872; // 90
        'h05b: dout <=  'sd1771; // 91
        'h05c: dout <=  'sd771; // 92
        'h05d: dout <=  'sd820; // 93
        'h05e: dout <=  'sd1570; // 94
        'h05f: dout <=  'sd1605; // 95
        'h060: dout <= -'sd816; // 96
        'h061: dout <=  'sd224; // 97
        'h062: dout <= -'sd2131; // 98
        'h063: dout <= -'sd260; // 99
        'h064: dout <=  'sd135; // 100
        'h065: dout <=  'sd243; // 101
        'h066: dout <= -'sd24; // 102
        'h067: dout <=  'sd124; // 103
        'h068: dout <=  'sd132; // 104
        'h069: dout <=  'sd2019; // 105
        'h06a: dout <= -'sd1000; // 106
        'h06b: dout <= -'sd1061; // 107
        'h06c: dout <= -'sd2025; // 108
        'h06d: dout <= -'sd1666; // 109
        'h06e: dout <= -'sd975; // 110
        'h06f: dout <= -'sd1519; // 111
        'h070: dout <= -'sd1948; // 112
        'h071: dout <= -'sd1380; // 113
        'h072: dout <= -'sd2142; // 114
        'h073: dout <= -'sd1343; // 115
        'h074: dout <=  'sd822; // 116
        'h075: dout <= -'sd818; // 117
        'h076: dout <=  'sd444; // 118
        'h077: dout <= -'sd1363; // 119
        'h078: dout <=  'sd1254; // 120
        'h079: dout <= -'sd611; // 121
        'h07a: dout <= -'sd1334; // 122
        'h07b: dout <=  'sd984; // 123
        'h07c: dout <=  'sd1759; // 124
        'h07d: dout <= -'sd1922; // 125
        'h07e: dout <= -'sd2034; // 126
        'h07f: dout <=  'sd426; // 127
        'h080: dout <= -'sd1589; // 128
        'h081: dout <=  'sd1420; // 129
        'h082: dout <= -'sd1588; // 130
        'h083: dout <=  'sd607; // 131
        'h084: dout <=  'sd852; // 132
        'h085: dout <= -'sd425; // 133
        'h086: dout <= -'sd1124; // 134
        'h087: dout <= -'sd419; // 135
        'h088: dout <=  'sd1818; // 136
        'h089: dout <=  'sd1514; // 137
        'h08a: dout <= -'sd1420; // 138
        'h08b: dout <=  'sd460; // 139
        'h08c: dout <= -'sd1417; // 140
        'h08d: dout <=  'sd606; // 141
        'h08e: dout <= -'sd1587; // 142
        'h08f: dout <= -'sd2032; // 143
        'h090: dout <=  'sd967; // 144
        'h091: dout <= -'sd1699; // 145
        'h092: dout <=  'sd1047; // 146
        'h093: dout <=  'sd382; // 147
        'h094: dout <= -'sd255; // 148
        'h095: dout <= -'sd1941; // 149
        'h096: dout <=  'sd1130; // 150
        'h097: dout <= -'sd553; // 151
        'h098: dout <=  'sd1996; // 152
        'h099: dout <=  'sd1003; // 153
        'h09a: dout <=  'sd811; // 154
        'h09b: dout <=  'sd1506; // 155
        'h09c: dout <= -'sd887; // 156
        'h09d: dout <=  'sd549; // 157
        'h09e: dout <=  'sd764; // 158
        'h09f: dout <=  'sd2175; // 159
        'h0a0: dout <= -'sd2243; // 160
        'h0a1: dout <= -'sd1278; // 161
        'h0a2: dout <= -'sd1278; // 162
        'h0a3: dout <= -'sd119; // 163
        'h0a4: dout <=  'sd1819; // 164
        'h0a5: dout <=  'sd1855; // 165
        'h0a6: dout <= -'sd2193; // 166
        'h0a7: dout <= -'sd1352; // 167
        'h0a8: dout <= -'sd1595; // 168
        'h0a9: dout <= -'sd1341; // 169
        'h0aa: dout <=  'sd1716; // 170
        'h0ab: dout <= -'sd840; // 171
        'h0ac: dout <= -'sd422; // 172
        'h0ad: dout <= -'sd107; // 173
        'h0ae: dout <=  'sd704; // 174
        'h0af: dout <= -'sd785; // 175
        'h0b0: dout <=  'sd233; // 176
        'h0b1: dout <=  'sd2214; // 177
        'h0b2: dout <=  'sd1927; // 178
        'h0b3: dout <=  'sd525; // 179
        'h0b4: dout <= -'sd458; // 180
        'h0b5: dout <= -'sd754; // 181
        'h0b6: dout <= -'sd2055; // 182
        'h0b7: dout <= -'sd1807; // 183
        'h0b8: dout <=  'sd1116; // 184
        'h0b9: dout <=  'sd424; // 185
        'h0ba: dout <= -'sd77; // 186
        'h0bb: dout <= -'sd1330; // 187
        'h0bc: dout <= -'sd468; // 188
        'h0bd: dout <=  'sd1642; // 189
        'h0be: dout <=  'sd627; // 190
        'h0bf: dout <=  'sd1710; // 191
        'h0c0: dout <=  'sd2027; // 192
        'h0c1: dout <= -'sd1138; // 193
        'h0c2: dout <= -'sd548; // 194
        'h0c3: dout <= -'sd2077; // 195
        'h0c4: dout <= -'sd1611; // 196
        'h0c5: dout <= -'sd1965; // 197
        'h0c6: dout <= -'sd799; // 198
        'h0c7: dout <=  'sd271; // 199
        'h0c8: dout <=  'sd2190; // 200
        'h0c9: dout <=  'sd1983; // 201
        'h0ca: dout <= -'sd234; // 202
        'h0cb: dout <= -'sd180; // 203
        'h0cc: dout <= -'sd628; // 204
        'h0cd: dout <=  'sd90; // 205
        'h0ce: dout <= -'sd954; // 206
        'h0cf: dout <=  'sd209; // 207
        'h0d0: dout <=  'sd1515; // 208
        'h0d1: dout <= -'sd993; // 209
        'h0d2: dout <=  'sd27; // 210
        'h0d3: dout <= -'sd97; // 211
        'h0d4: dout <= -'sd349; // 212
        'h0d5: dout <=  'sd2132; // 213
        'h0d6: dout <= -'sd417; // 214
        'h0d7: dout <= -'sd313; // 215
        'h0d8: dout <=  'sd1153; // 216
        'h0d9: dout <= -'sd1564; // 217
        'h0da: dout <=  'sd869; // 218
        'h0db: dout <= -'sd1634; // 219
        'h0dc: dout <= -'sd2049; // 220
        'h0dd: dout <= -'sd2206; // 221
        'h0de: dout <=  'sd1491; // 222
        'h0df: dout <=  'sd1831; // 223
        'h0e0: dout <= -'sd16; // 224
        'h0e1: dout <=  'sd1690; // 225
        'h0e2: dout <=  'sd2252; // 226
        'h0e3: dout <=  'sd1987; // 227
        'h0e4: dout <=  'sd1077; // 228
        'h0e5: dout <=  'sd1207; // 229
        'h0e6: dout <=  'sd699; // 230
        'h0e7: dout <= -'sd23; // 231
        'h0e8: dout <=  'sd1534; // 232
        'h0e9: dout <= -'sd1202; // 233
        'h0ea: dout <= -'sd38; // 234
        'h0eb: dout <=  'sd198; // 235
        'h0ec: dout <=  'sd296; // 236
        'h0ed: dout <=  'sd827; // 237
        'h0ee: dout <= -'sd1320; // 238
        'h0ef: dout <=  'sd1856; // 239
        'h0f0: dout <= -'sd1802; // 240
        'h0f1: dout <=  'sd769; // 241
        'h0f2: dout <=  'sd1806; // 242
        'h0f3: dout <= -'sd1595; // 243
        'h0f4: dout <= -'sd834; // 244
        'h0f5: dout <=  'sd1025; // 245
        'h0f6: dout <=  'sd556; // 246
        'h0f7: dout <= -'sd1585; // 247
        'h0f8: dout <=  'sd464; // 248
        'h0f9: dout <= -'sd1564; // 249
        'h0fa: dout <= -'sd132; // 250
        'h0fb: dout <= -'sd2197; // 251
        'h0fc: dout <= -'sd296; // 252
        'h0fd: dout <= -'sd798; // 253
        'h0fe: dout <=  'sd626; // 254
        'h0ff: dout <=  'sd903; // 255
        'h100: dout <=  'sd2080; // 256
        'h101: dout <=  'sd22; // 257
        'h102: dout <=  'sd1856; // 258
        'h103: dout <= -'sd792; // 259
        'h104: dout <= -'sd941; // 260
        'h105: dout <= -'sd1016; // 261
        'h106: dout <= -'sd103; // 262
        'h107: dout <=  'sd1092; // 263
        'h108: dout <= -'sd1917; // 264
        'h109: dout <= -'sd1743; // 265
        'h10a: dout <= -'sd175; // 266
        'h10b: dout <=  'sd1032; // 267
        'h10c: dout <=  'sd708; // 268
        'h10d: dout <=  'sd117; // 269
        'h10e: dout <=  'sd1380; // 270
        'h10f: dout <= -'sd650; // 271
        'h110: dout <= -'sd1519; // 272
        'h111: dout <=  'sd114; // 273
        'h112: dout <=  'sd1510; // 274
        'h113: dout <=  'sd1978; // 275
        'h114: dout <=  'sd1642; // 276
        'h115: dout <= -'sd27; // 277
        'h116: dout <=  'sd846; // 278
        'h117: dout <= -'sd873; // 279
        'h118: dout <=  'sd242; // 280
        'h119: dout <=  'sd597; // 281
        'h11a: dout <= -'sd1038; // 282
        'h11b: dout <=  'sd2110; // 283
        'h11c: dout <=  'sd699; // 284
        'h11d: dout <=  'sd78; // 285
        'h11e: dout <= -'sd92; // 286
        'h11f: dout <=  'sd1652; // 287
        'h120: dout <= -'sd442; // 288
        'h121: dout <= -'sd1656; // 289
        'h122: dout <= -'sd838; // 290
        'h123: dout <=  'sd1635; // 291
        'h124: dout <= -'sd330; // 292
        'h125: dout <= -'sd2236; // 293
        'h126: dout <=  'sd1819; // 294
        'h127: dout <=  'sd1384; // 295
        'h128: dout <=  'sd248; // 296
        'h129: dout <= -'sd1063; // 297
        'h12a: dout <= -'sd963; // 298
        'h12b: dout <= -'sd1040; // 299
        'h12c: dout <= -'sd1135; // 300
        'h12d: dout <=  'sd230; // 301
        'h12e: dout <= -'sd2286; // 302
        'h12f: dout <= -'sd988; // 303
        'h130: dout <= -'sd2001; // 304
        'h131: dout <= -'sd902; // 305
        'h132: dout <=  'sd1379; // 306
        'h133: dout <= -'sd1747; // 307
        'h134: dout <=  'sd626; // 308
        'h135: dout <= -'sd1632; // 309
        'h136: dout <=  'sd104; // 310
        'h137: dout <=  'sd1475; // 311
        'h138: dout <= -'sd1503; // 312
        'h139: dout <=  'sd1793; // 313
        'h13a: dout <=  'sd315; // 314
        'h13b: dout <= -'sd886; // 315
        'h13c: dout <= -'sd381; // 316
        'h13d: dout <= -'sd2190; // 317
        'h13e: dout <=  'sd829; // 318
        'h13f: dout <= -'sd53; // 319
        'h140: dout <= -'sd1352; // 320
        'h141: dout <=  'sd754; // 321
        'h142: dout <= -'sd291; // 322
        'h143: dout <=  'sd956; // 323
        'h144: dout <=  'sd990; // 324
        'h145: dout <=  'sd883; // 325
        'h146: dout <=  'sd623; // 326
        'h147: dout <= -'sd141; // 327
        'h148: dout <= -'sd914; // 328
        'h149: dout <=  'sd548; // 329
        'h14a: dout <=  'sd1514; // 330
        'h14b: dout <= -'sd341; // 331
        'h14c: dout <= -'sd1909; // 332
        'h14d: dout <=  'sd667; // 333
        'h14e: dout <=  'sd682; // 334
        'h14f: dout <= -'sd1192; // 335
        'h150: dout <= -'sd1846; // 336
        'h151: dout <=  'sd2120; // 337
        'h152: dout <= -'sd1971; // 338
        'h153: dout <=  'sd2022; // 339
        'h154: dout <= -'sd1768; // 340
        'h155: dout <=  'sd213; // 341
        'h156: dout <=  'sd1896; // 342
        'h157: dout <=  'sd2111; // 343
        'h158: dout <= -'sd1722; // 344
        'h159: dout <= -'sd819; // 345
        'h15a: dout <=  'sd190; // 346
        'h15b: dout <=  'sd1273; // 347
        'h15c: dout <= -'sd596; // 348
        'h15d: dout <= -'sd1523; // 349
        'h15e: dout <=  'sd966; // 350
        'h15f: dout <=  'sd892; // 351
        'h160: dout <= -'sd1788; // 352
        'h161: dout <=  'sd1223; // 353
        'h162: dout <= -'sd240; // 354
        'h163: dout <=  'sd1754; // 355
        'h164: dout <=  'sd2183; // 356
        'h165: dout <=  'sd190; // 357
        'h166: dout <=  'sd438; // 358
        'h167: dout <=  'sd1981; // 359
        'h168: dout <=  'sd1266; // 360
        'h169: dout <= -'sd233; // 361
        'h16a: dout <= -'sd117; // 362
        'h16b: dout <=  'sd1684; // 363
        'h16c: dout <= -'sd1948; // 364
        'h16d: dout <= -'sd1630; // 365
        'h16e: dout <= -'sd2074; // 366
        'h16f: dout <= -'sd1131; // 367
        'h170: dout <=  'sd1648; // 368
        'h171: dout <= -'sd749; // 369
        'h172: dout <=  'sd1417; // 370
        'h173: dout <= -'sd2172; // 371
        'h174: dout <= -'sd1111; // 372
        'h175: dout <= -'sd2088; // 373
        'h176: dout <= -'sd2121; // 374
        'h177: dout <=  'sd415; // 375
        'h178: dout <= -'sd366; // 376
        'h179: dout <=  'sd394; // 377
        'h17a: dout <=  'sd2002; // 378
        'h17b: dout <= -'sd1498; // 379
        'h17c: dout <= -'sd1634; // 380
        'h17d: dout <=  'sd987; // 381
        'h17e: dout <= -'sd1567; // 382
        'h17f: dout <= -'sd1064; // 383
        'h180: dout <= -'sd1117; // 384
        'h181: dout <= -'sd1147; // 385
        'h182: dout <=  'sd1484; // 386
        'h183: dout <= -'sd50; // 387
        'h184: dout <=  'sd709; // 388
        'h185: dout <= -'sd758; // 389
        'h186: dout <= -'sd2162; // 390
        'h187: dout <=  'sd2249; // 391
        'h188: dout <=  'sd2166; // 392
        'h189: dout <=  'sd101; // 393
        'h18a: dout <=  'sd1048; // 394
        'h18b: dout <=  'sd2249; // 395
        'h18c: dout <=  'sd855; // 396
        'h18d: dout <= -'sd1773; // 397
        'h18e: dout <=  'sd255; // 398
        'h18f: dout <= -'sd413; // 399
        'h190: dout <=  'sd1205; // 400
        'h191: dout <=  'sd261; // 401
        'h192: dout <=  'sd1321; // 402
        'h193: dout <= -'sd216; // 403
        'h194: dout <= -'sd1397; // 404
        'h195: dout <= -'sd285; // 405
        'h196: dout <= -'sd362; // 406
        'h197: dout <=  'sd1654; // 407
        'h198: dout <=  'sd158; // 408
        'h199: dout <=  'sd1951; // 409
        'h19a: dout <=  'sd2222; // 410
        'h19b: dout <= -'sd455; // 411
        'h19c: dout <= -'sd1565; // 412
        'h19d: dout <= -'sd1751; // 413
        'h19e: dout <= -'sd1541; // 414
        'h19f: dout <=  'sd1164; // 415
        'h1a0: dout <= -'sd352; // 416
        'h1a1: dout <=  'sd1731; // 417
        'h1a2: dout <= -'sd243; // 418
        'h1a3: dout <= -'sd2100; // 419
        'h1a4: dout <=  'sd121; // 420
        'h1a5: dout <=  'sd1714; // 421
        'h1a6: dout <= -'sd84; // 422
        'h1a7: dout <=  'sd528; // 423
        'h1a8: dout <=  'sd2135; // 424
        'h1a9: dout <=  'sd1250; // 425
        'h1aa: dout <= -'sd746; // 426
        'h1ab: dout <= -'sd86; // 427
        'h1ac: dout <= -'sd8; // 428
        'h1ad: dout <=  'sd1993; // 429
        'h1ae: dout <= -'sd2007; // 430
        'h1af: dout <=  'sd2110; // 431
        'h1b0: dout <= -'sd1136; // 432
        'h1b1: dout <= -'sd249; // 433
        'h1b2: dout <= -'sd814; // 434
        'h1b3: dout <= -'sd693; // 435
        'h1b4: dout <=  'sd1300; // 436
        'h1b5: dout <=  'sd563; // 437
        'h1b6: dout <= -'sd45; // 438
        'h1b7: dout <=  'sd299; // 439
        'h1b8: dout <=  'sd1709; // 440
        'h1b9: dout <= -'sd1643; // 441
        'h1ba: dout <= -'sd427; // 442
        'h1bb: dout <=  'sd113; // 443
        'h1bc: dout <=  'sd1975; // 444
        'h1bd: dout <=  'sd2075; // 445
        'h1be: dout <=  'sd742; // 446
        'h1bf: dout <=  'sd1671; // 447
        'h1c0: dout <= -'sd1368; // 448
        'h1c1: dout <= -'sd2142; // 449
        'h1c2: dout <=  'sd349; // 450
        'h1c3: dout <= -'sd275; // 451
        'h1c4: dout <=  'sd359; // 452
        'h1c5: dout <=  'sd1415; // 453
        'h1c6: dout <=  'sd752; // 454
        'h1c7: dout <=  'sd1639; // 455
        'h1c8: dout <=  'sd1518; // 456
        'h1c9: dout <= -'sd1561; // 457
        'h1ca: dout <=  'sd891; // 458
        'h1cb: dout <= -'sd2223; // 459
        'h1cc: dout <=  'sd602; // 460
        'h1cd: dout <=  'sd1042; // 461
        'h1ce: dout <= -'sd988; // 462
        'h1cf: dout <= -'sd445; // 463
        'h1d0: dout <=  'sd240; // 464
        'h1d1: dout <= -'sd1589; // 465
        'h1d2: dout <=  'sd2151; // 466
        'h1d3: dout <= -'sd218; // 467
        'h1d4: dout <= -'sd1358; // 468
        'h1d5: dout <= -'sd975; // 469
        'h1d6: dout <=  'sd1533; // 470
        'h1d7: dout <=  'sd2254; // 471
        'h1d8: dout <= -'sd1062; // 472
        'h1d9: dout <=  'sd1580; // 473
        'h1da: dout <= -'sd2292; // 474
        'h1db: dout <=  'sd428; // 475
        'h1dc: dout <= -'sd1313; // 476
        'h1dd: dout <=  'sd1214; // 477
        'h1de: dout <= -'sd645; // 478
        'h1df: dout <=  'sd460; // 479
        'h1e0: dout <= -'sd1555; // 480
        'h1e1: dout <= -'sd1357; // 481
        'h1e2: dout <=  'sd861; // 482
        'h1e3: dout <=  'sd445; // 483
        'h1e4: dout <= -'sd1796; // 484
        'h1e5: dout <= -'sd1927; // 485
        'h1e6: dout <=  'sd776; // 486
        'h1e7: dout <=  'sd437; // 487
        'h1e8: dout <=  'sd1754; // 488
        'h1e9: dout <= -'sd163; // 489
        'h1ea: dout <= -'sd1154; // 490
        'h1eb: dout <= -'sd1813; // 491
        'h1ec: dout <=  'sd1041; // 492
        'h1ed: dout <= -'sd2246; // 493
        'h1ee: dout <=  'sd1788; // 494
        'h1ef: dout <=  'sd736; // 495
        'h1f0: dout <= -'sd1931; // 496
        'h1f1: dout <= -'sd2245; // 497
        'h1f2: dout <= -'sd751; // 498
        'h1f3: dout <= -'sd79; // 499
        'h1f4: dout <= -'sd698; // 500
        'h1f5: dout <=  'sd878; // 501
        'h1f6: dout <=  'sd239; // 502
        'h1f7: dout <=  'sd2206; // 503
        'h1f8: dout <=  'sd947; // 504
        'h1f9: dout <= -'sd1998; // 505
        'h1fa: dout <= -'sd371; // 506
        'h1fb: dout <=  'sd547; // 507
        'h1fc: dout <= -'sd448; // 508
        'h1fd: dout <=  'sd1217; // 509
        'h1fe: dout <=  'sd71; // 510
        'h1ff: dout <= -'sd247; // 511
        'h200: dout <= -'sd1995; // 512
        'h201: dout <=  'sd20; // 513
        'h202: dout <=  'sd2139; // 514
        'h203: dout <=  'sd784; // 515
        'h204: dout <=  'sd2075; // 516
        'h205: dout <=  'sd1747; // 517
        'h206: dout <= -'sd1212; // 518
        'h207: dout <=  'sd1264; // 519
        'h208: dout <=  'sd488; // 520
        'h209: dout <=  'sd1002; // 521
        'h20a: dout <=  'sd1676; // 522
        'h20b: dout <= -'sd1652; // 523
        'h20c: dout <= -'sd1988; // 524
        'h20d: dout <=  'sd1710; // 525
        'h20e: dout <=  'sd843; // 526
        'h20f: dout <= -'sd1718; // 527
        'h210: dout <= -'sd1957; // 528
        'h211: dout <= -'sd361; // 529
        'h212: dout <=  'sd791; // 530
        'h213: dout <= -'sd1461; // 531
        'h214: dout <=  'sd2034; // 532
        'h215: dout <= -'sd1470; // 533
        'h216: dout <= -'sd282; // 534
        'h217: dout <= -'sd1455; // 535
        'h218: dout <=  'sd1365; // 536
        'h219: dout <=  'sd2268; // 537
        'h21a: dout <=  'sd1679; // 538
        'h21b: dout <=  'sd1782; // 539
        'h21c: dout <=  'sd1788; // 540
        'h21d: dout <= -'sd1524; // 541
        'h21e: dout <=  'sd894; // 542
        'h21f: dout <=  'sd663; // 543
        'h220: dout <=  'sd2187; // 544
        'h221: dout <= -'sd196; // 545
        'h222: dout <= -'sd199; // 546
        'h223: dout <=  'sd860; // 547
        'h224: dout <=  'sd766; // 548
        'h225: dout <= -'sd2105; // 549
        'h226: dout <= -'sd2157; // 550
        'h227: dout <= -'sd2123; // 551
        'h228: dout <= -'sd482; // 552
        'h229: dout <=  'sd1165; // 553
        'h22a: dout <=  'sd1174; // 554
        'h22b: dout <= -'sd1990; // 555
        'h22c: dout <= -'sd1097; // 556
        'h22d: dout <=  'sd1994; // 557
        'h22e: dout <= -'sd922; // 558
        'h22f: dout <= -'sd903; // 559
        'h230: dout <= -'sd330; // 560
        'h231: dout <= -'sd2156; // 561
        'h232: dout <= -'sd692; // 562
        'h233: dout <=  'sd505; // 563
        'h234: dout <=  'sd254; // 564
        'h235: dout <= -'sd1907; // 565
        'h236: dout <=  'sd1079; // 566
        'h237: dout <= -'sd485; // 567
        'h238: dout <=  'sd2245; // 568
        'h239: dout <=  'sd1027; // 569
        'h23a: dout <= -'sd424; // 570
        'h23b: dout <=  'sd255; // 571
        'h23c: dout <=  'sd87; // 572
        'h23d: dout <=  'sd752; // 573
        'h23e: dout <= -'sd287; // 574
        'h23f: dout <=  'sd2068; // 575
        'h240: dout <= -'sd1636; // 576
        'h241: dout <= -'sd33; // 577
        'h242: dout <= -'sd344; // 578
        'h243: dout <=  'sd247; // 579
        'h244: dout <= -'sd170; // 580
        'h245: dout <= -'sd674; // 581
        'h246: dout <= -'sd2026; // 582
        'h247: dout <= -'sd960; // 583
        'h248: dout <= -'sd1927; // 584
        'h249: dout <= -'sd2024; // 585
        'h24a: dout <= -'sd1614; // 586
        'h24b: dout <= -'sd764; // 587
        'h24c: dout <= -'sd2188; // 588
        'h24d: dout <= -'sd1868; // 589
        'h24e: dout <=  'sd602; // 590
        'h24f: dout <= -'sd373; // 591
        'h250: dout <= -'sd249; // 592
        'h251: dout <=  'sd620; // 593
        'h252: dout <=  'sd1996; // 594
        'h253: dout <=  'sd1621; // 595
        'h254: dout <=  'sd1094; // 596
        'h255: dout <=  'sd1658; // 597
        'h256: dout <=  'sd2221; // 598
        'h257: dout <=  'sd983; // 599
        'h258: dout <= -'sd1256; // 600
        'h259: dout <= -'sd2072; // 601
        'h25a: dout <=  'sd2005; // 602
        'h25b: dout <= -'sd562; // 603
        'h25c: dout <= -'sd1045; // 604
        'h25d: dout <= -'sd1246; // 605
        'h25e: dout <=  'sd1922; // 606
        'h25f: dout <=  'sd15; // 607
        'h260: dout <= -'sd783; // 608
        'h261: dout <=  'sd876; // 609
        'h262: dout <= -'sd952; // 610
        'h263: dout <=  'sd2042; // 611
        'h264: dout <=  'sd1515; // 612
        'h265: dout <=  'sd1122; // 613
        'h266: dout <=  'sd785; // 614
        'h267: dout <=  'sd1414; // 615
        'h268: dout <= -'sd442; // 616
        'h269: dout <= -'sd1450; // 617
        'h26a: dout <=  'sd2142; // 618
        'h26b: dout <=  'sd32; // 619
        'h26c: dout <=  'sd2290; // 620
        'h26d: dout <=  'sd1141; // 621
        'h26e: dout <=  'sd614; // 622
        'h26f: dout <=  'sd1059; // 623
        'h270: dout <= -'sd877; // 624
        'h271: dout <=  'sd757; // 625
        'h272: dout <= -'sd2074; // 626
        'h273: dout <=  'sd806; // 627
        'h274: dout <= -'sd1963; // 628
        'h275: dout <= -'sd1619; // 629
        'h276: dout <=  'sd1263; // 630
        'h277: dout <= -'sd1448; // 631
        'h278: dout <= -'sd518; // 632
        'h279: dout <= -'sd2157; // 633
        'h27a: dout <= -'sd481; // 634
        'h27b: dout <= -'sd348; // 635
        'h27c: dout <=  'sd70; // 636
        'h27d: dout <=  'sd543; // 637
        'h27e: dout <= -'sd1116; // 638
        'h27f: dout <=  'sd1601; // 639
        'h280: dout <= -'sd130; // 640
        'h281: dout <=  'sd686; // 641
        'h282: dout <=  'sd336; // 642
        'h283: dout <=  'sd1306; // 643
        'h284: dout <=  'sd1945; // 644
        'h285: dout <= -'sd743; // 645
        'h286: dout <=  'sd1829; // 646
        'h287: dout <=  'sd214; // 647
        'h288: dout <=  'sd1255; // 648
        'h289: dout <=  'sd754; // 649
        'h28a: dout <=  'sd422; // 650
        'h28b: dout <= -'sd867; // 651
        'h28c: dout <=  'sd2165; // 652
        'h28d: dout <= -'sd403; // 653
        'h28e: dout <= -'sd1336; // 654
        'h28f: dout <= -'sd428; // 655
        'h290: dout <=  'sd755; // 656
        'h291: dout <= -'sd158; // 657
        'h292: dout <= -'sd10; // 658
        'h293: dout <=  'sd1417; // 659
        'h294: dout <=  'sd210; // 660
        'h295: dout <= -'sd1668; // 661
        'h296: dout <=  'sd2153; // 662
        'h297: dout <= -'sd625; // 663
        'h298: dout <= -'sd2291; // 664
        'h299: dout <=  'sd131; // 665
        'h29a: dout <= -'sd1081; // 666
        'h29b: dout <= -'sd369; // 667
        'h29c: dout <=  'sd714; // 668
        'h29d: dout <= -'sd1271; // 669
        'h29e: dout <=  'sd62; // 670
        'h29f: dout <=  'sd1542; // 671
        'h2a0: dout <=  'sd2025; // 672
        'h2a1: dout <= -'sd672; // 673
        'h2a2: dout <=  'sd1066; // 674
        'h2a3: dout <=  'sd901; // 675
        'h2a4: dout <=  'sd546; // 676
        'h2a5: dout <= -'sd76; // 677
        'h2a6: dout <= -'sd358; // 678
        'h2a7: dout <= -'sd841; // 679
        'h2a8: dout <=  'sd263; // 680
        'h2a9: dout <= -'sd1130; // 681
        'h2aa: dout <=  'sd1234; // 682
        'h2ab: dout <=  'sd1171; // 683
        'h2ac: dout <= -'sd1617; // 684
        'h2ad: dout <=  'sd1042; // 685
        'h2ae: dout <=  'sd627; // 686
        'h2af: dout <= -'sd27; // 687
        'h2b0: dout <=  'sd1603; // 688
        'h2b1: dout <=  'sd1107; // 689
        'h2b2: dout <= -'sd1628; // 690
        'h2b3: dout <=  'sd42; // 691
        'h2b4: dout <= -'sd706; // 692
        'h2b5: dout <= -'sd888; // 693
        'h2b6: dout <=  'sd513; // 694
        'h2b7: dout <= -'sd580; // 695
        'h2b8: dout <= -'sd511; // 696
        'h2b9: dout <=  'sd147; // 697
        'h2ba: dout <= -'sd1741; // 698
        'h2bb: dout <= -'sd586; // 699
        'h2bc: dout <=  'sd229; // 700
        'h2bd: dout <= -'sd94; // 701
        'h2be: dout <= -'sd1673; // 702
        'h2bf: dout <=  'sd87; // 703
        'h2c0: dout <= -'sd463; // 704
        'h2c1: dout <= -'sd1178; // 705
        'h2c2: dout <= -'sd179; // 706
        'h2c3: dout <=  'sd1755; // 707
        'h2c4: dout <=  'sd1826; // 708
        'h2c5: dout <=  'sd1317; // 709
        'h2c6: dout <= -'sd1325; // 710
        'h2c7: dout <= -'sd407; // 711
        'h2c8: dout <= -'sd2236; // 712
        'h2c9: dout <=  'sd967; // 713
        'h2ca: dout <= -'sd2176; // 714
        'h2cb: dout <=  'sd1652; // 715
        'h2cc: dout <=  'sd1765; // 716
        'h2cd: dout <=  'sd525; // 717
        'h2ce: dout <=  'sd1670; // 718
        'h2cf: dout <=  'sd285; // 719
        'h2d0: dout <=  'sd1968; // 720
        'h2d1: dout <=  'sd322; // 721
        'h2d2: dout <=  'sd427; // 722
        'h2d3: dout <=  'sd1799; // 723
        'h2d4: dout <=  'sd1712; // 724
        'h2d5: dout <= -'sd276; // 725
        'h2d6: dout <= -'sd1238; // 726
        'h2d7: dout <=  'sd930; // 727
        'h2d8: dout <= -'sd498; // 728
        'h2d9: dout <=  'sd1446; // 729
        'h2da: dout <= -'sd1244; // 730
        'h2db: dout <= -'sd249; // 731
        'h2dc: dout <= -'sd1567; // 732
        'h2dd: dout <=  'sd1587; // 733
        'h2de: dout <=  'sd331; // 734
        'h2df: dout <=  'sd1911; // 735
        'h2e0: dout <= -'sd2238; // 736
        'h2e1: dout <= -'sd1693; // 737
        'h2e2: dout <=  'sd381; // 738
        'h2e3: dout <=  'sd981; // 739
        'h2e4: dout <=  'sd1114; // 740
        'h2e5: dout <=  'sd805; // 741
        'h2e6: dout <= -'sd98; // 742
        'h2e7: dout <=  'sd781; // 743
        'h2e8: dout <= -'sd239; // 744
        'h2e9: dout <=  'sd1909; // 745
        'h2ea: dout <=  'sd2227; // 746
        'h2eb: dout <=  'sd69; // 747
        'h2ec: dout <= -'sd1235; // 748
        'h2ed: dout <= -'sd1286; // 749
        'h2ee: dout <=  'sd19; // 750
        'h2ef: dout <= -'sd468; // 751
        'h2f0: dout <=  'sd640; // 752
        'h2f1: dout <= -'sd1705; // 753
        'h2f2: dout <=  'sd348; // 754
        'h2f3: dout <=  'sd1790; // 755
        'h2f4: dout <= -'sd1415; // 756
        'h2f5: dout <=  'sd2144; // 757
        'h2f6: dout <=  'sd1890; // 758
        'h2f7: dout <= -'sd1477; // 759
        'h2f8: dout <=  'sd591; // 760
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hq1_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <=  'sd52177; // 0
        'h001: dout <= -'sd10255; // 1
        'h002: dout <= -'sd7800; // 2
        'h003: dout <=  'sd54944; // 3
        'h004: dout <= -'sd50265; // 4
        'h005: dout <= -'sd14159; // 5
        'h006: dout <=  'sd17307; // 6
        'h007: dout <=  'sd32823; // 7
        'h008: dout <=  'sd46203; // 8
        'h009: dout <=  'sd3771; // 9
        'h00a: dout <= -'sd41573; // 10
        'h00b: dout <= -'sd54916; // 11
        'h00c: dout <= -'sd48040; // 12
        'h00d: dout <=  'sd15636; // 13
        'h00e: dout <= -'sd37342; // 14
        'h00f: dout <=  'sd29429; // 15
        'h010: dout <= -'sd24222; // 16
        'h011: dout <= -'sd44803; // 17
        'h012: dout <=  'sd43418; // 18
        'h013: dout <=  'sd11365; // 19
        'h014: dout <= -'sd56619; // 20
        'h015: dout <=  'sd42265; // 21
        'h016: dout <=  'sd43227; // 22
        'h017: dout <= -'sd18487; // 23
        'h018: dout <=  'sd6837; // 24
        'h019: dout <= -'sd46253; // 25
        'h01a: dout <=  'sd12117; // 26
        'h01b: dout <=  'sd43260; // 27
        'h01c: dout <=  'sd14749; // 28
        'h01d: dout <=  'sd43866; // 29
        'h01e: dout <= -'sd56890; // 30
        'h01f: dout <=  'sd35721; // 31
        'h020: dout <=  'sd39671; // 32
        'h021: dout <= -'sd10652; // 33
        'h022: dout <= -'sd6809; // 34
        'h023: dout <=  'sd2036; // 35
        'h024: dout <=  'sd30307; // 36
        'h025: dout <=  'sd27541; // 37
        'h026: dout <= -'sd24658; // 38
        'h027: dout <=  'sd2717; // 39
        'h028: dout <= -'sd51417; // 40
        'h029: dout <= -'sd2296; // 41
        'h02a: dout <= -'sd18127; // 42
        'h02b: dout <=  'sd11372; // 43
        'h02c: dout <=  'sd29440; // 44
        'h02d: dout <= -'sd32253; // 45
        'h02e: dout <= -'sd31109; // 46
        'h02f: dout <= -'sd19945; // 47
        'h030: dout <=  'sd52786; // 48
        'h031: dout <= -'sd15810; // 49
        'h032: dout <=  'sd16882; // 50
        'h033: dout <=  'sd30758; // 51
        'h034: dout <= -'sd47681; // 52
        'h035: dout <= -'sd12309; // 53
        'h036: dout <=  'sd56866; // 54
        'h037: dout <=  'sd42867; // 55
        'h038: dout <= -'sd28568; // 56
        'h039: dout <=  'sd10695; // 57
        'h03a: dout <= -'sd17021; // 58
        'h03b: dout <= -'sd30303; // 59
        'h03c: dout <= -'sd44632; // 60
        'h03d: dout <=  'sd44278; // 61
        'h03e: dout <= -'sd48471; // 62
        'h03f: dout <= -'sd56867; // 63
        'h040: dout <=  'sd10991; // 64
        'h041: dout <=  'sd15525; // 65
        'h042: dout <=  'sd11310; // 66
        'h043: dout <=  'sd47824; // 67
        'h044: dout <=  'sd15941; // 68
        'h045: dout <= -'sd20444; // 69
        'h046: dout <= -'sd48231; // 70
        'h047: dout <= -'sd8374; // 71
        'h048: dout <=  'sd2908; // 72
        'h049: dout <=  'sd21365; // 73
        'h04a: dout <= -'sd27110; // 74
        'h04b: dout <=  'sd3002; // 75
        'h04c: dout <= -'sd37728; // 76
        'h04d: dout <=  'sd27403; // 77
        'h04e: dout <= -'sd46481; // 78
        'h04f: dout <=  'sd40174; // 79
        'h050: dout <=  'sd15371; // 80
        'h051: dout <=  'sd13028; // 81
        'h052: dout <=  'sd21341; // 82
        'h053: dout <= -'sd50704; // 83
        'h054: dout <=  'sd43810; // 84
        'h055: dout <= -'sd28279; // 85
        'h056: dout <=  'sd21343; // 86
        'h057: dout <= -'sd54150; // 87
        'h058: dout <=  'sd8643; // 88
        'h059: dout <= -'sd19130; // 89
        'h05a: dout <= -'sd35691; // 90
        'h05b: dout <=  'sd9417; // 91
        'h05c: dout <=  'sd55473; // 92
        'h05d: dout <= -'sd7529; // 93
        'h05e: dout <=  'sd38411; // 94
        'h05f: dout <=  'sd4994; // 95
        'h060: dout <=  'sd42328; // 96
        'h061: dout <= -'sd39838; // 97
        'h062: dout <=  'sd26133; // 98
        'h063: dout <=  'sd1659; // 99
        'h064: dout <= -'sd40047; // 100
        'h065: dout <=  'sd53038; // 101
        'h066: dout <= -'sd46813; // 102
        'h067: dout <=  'sd28403; // 103
        'h068: dout <=  'sd44678; // 104
        'h069: dout <=  'sd54475; // 105
        'h06a: dout <= -'sd29319; // 106
        'h06b: dout <= -'sd51116; // 107
        'h06c: dout <= -'sd53564; // 108
        'h06d: dout <= -'sd2166; // 109
        'h06e: dout <=  'sd45639; // 110
        'h06f: dout <=  'sd3719; // 111
        'h070: dout <=  'sd42284; // 112
        'h071: dout <= -'sd45547; // 113
        'h072: dout <=  'sd19506; // 114
        'h073: dout <=  'sd33272; // 115
        'h074: dout <= -'sd8603; // 116
        'h075: dout <=  'sd42727; // 117
        'h076: dout <=  'sd10577; // 118
        'h077: dout <=  'sd19384; // 119
        'h078: dout <= -'sd15999; // 120
        'h079: dout <= -'sd27987; // 121
        'h07a: dout <=  'sd13658; // 122
        'h07b: dout <= -'sd50381; // 123
        'h07c: dout <=  'sd27792; // 124
        'h07d: dout <=  'sd21228; // 125
        'h07e: dout <=  'sd56486; // 126
        'h07f: dout <= -'sd36427; // 127
        'h080: dout <= -'sd35573; // 128
        'h081: dout <=  'sd12203; // 129
        'h082: dout <=  'sd21423; // 130
        'h083: dout <=  'sd10169; // 131
        'h084: dout <= -'sd34229; // 132
        'h085: dout <= -'sd44760; // 133
        'h086: dout <=  'sd20951; // 134
        'h087: dout <=  'sd4149; // 135
        'h088: dout <= -'sd31178; // 136
        'h089: dout <= -'sd25733; // 137
        'h08a: dout <=  'sd21107; // 138
        'h08b: dout <= -'sd28221; // 139
        'h08c: dout <=  'sd12562; // 140
        'h08d: dout <=  'sd2560; // 141
        'h08e: dout <= -'sd9089; // 142
        'h08f: dout <= -'sd2131; // 143
        'h090: dout <=  'sd5834; // 144
        'h091: dout <= -'sd56613; // 145
        'h092: dout <=  'sd16060; // 146
        'h093: dout <=  'sd12124; // 147
        'h094: dout <= -'sd14994; // 148
        'h095: dout <=  'sd24101; // 149
        'h096: dout <=  'sd55441; // 150
        'h097: dout <= -'sd52896; // 151
        'h098: dout <=  'sd37567; // 152
        'h099: dout <=  'sd42236; // 153
        'h09a: dout <= -'sd21509; // 154
        'h09b: dout <= -'sd5387; // 155
        'h09c: dout <=  'sd3602; // 156
        'h09d: dout <= -'sd30574; // 157
        'h09e: dout <= -'sd48266; // 158
        'h09f: dout <=  'sd51642; // 159
        'h0a0: dout <=  'sd17011; // 160
        'h0a1: dout <= -'sd43858; // 161
        'h0a2: dout <=  'sd45456; // 162
        'h0a3: dout <=  'sd25528; // 163
        'h0a4: dout <=  'sd5970; // 164
        'h0a5: dout <=  'sd55591; // 165
        'h0a6: dout <= -'sd19970; // 166
        'h0a7: dout <= -'sd34032; // 167
        'h0a8: dout <= -'sd34347; // 168
        'h0a9: dout <= -'sd29130; // 169
        'h0aa: dout <=  'sd751; // 170
        'h0ab: dout <= -'sd2945; // 171
        'h0ac: dout <=  'sd46161; // 172
        'h0ad: dout <= -'sd39177; // 173
        'h0ae: dout <=  'sd12077; // 174
        'h0af: dout <= -'sd17878; // 175
        'h0b0: dout <= -'sd16580; // 176
        'h0b1: dout <= -'sd11198; // 177
        'h0b2: dout <= -'sd5048; // 178
        'h0b3: dout <= -'sd12024; // 179
        'h0b4: dout <= -'sd39604; // 180
        'h0b5: dout <=  'sd4501; // 181
        'h0b6: dout <=  'sd36231; // 182
        'h0b7: dout <=  'sd52086; // 183
        'h0b8: dout <=  'sd6163; // 184
        'h0b9: dout <=  'sd34591; // 185
        'h0ba: dout <= -'sd40003; // 186
        'h0bb: dout <=  'sd15721; // 187
        'h0bc: dout <=  'sd49795; // 188
        'h0bd: dout <= -'sd33531; // 189
        'h0be: dout <=  'sd51766; // 190
        'h0bf: dout <=  'sd48030; // 191
        'h0c0: dout <= -'sd25121; // 192
        'h0c1: dout <=  'sd42035; // 193
        'h0c2: dout <= -'sd38510; // 194
        'h0c3: dout <=  'sd13519; // 195
        'h0c4: dout <= -'sd31323; // 196
        'h0c5: dout <=  'sd25278; // 197
        'h0c6: dout <=  'sd47860; // 198
        'h0c7: dout <=  'sd30517; // 199
        'h0c8: dout <= -'sd38946; // 200
        'h0c9: dout <= -'sd38310; // 201
        'h0ca: dout <= -'sd50106; // 202
        'h0cb: dout <= -'sd38684; // 203
        'h0cc: dout <=  'sd14128; // 204
        'h0cd: dout <= -'sd37833; // 205
        'h0ce: dout <= -'sd40731; // 206
        'h0cf: dout <=  'sd13468; // 207
        'h0d0: dout <=  'sd3542; // 208
        'h0d1: dout <=  'sd3615; // 209
        'h0d2: dout <=  'sd16455; // 210
        'h0d3: dout <= -'sd19475; // 211
        'h0d4: dout <=  'sd19218; // 212
        'h0d5: dout <=  'sd36820; // 213
        'h0d6: dout <= -'sd29556; // 214
        'h0d7: dout <= -'sd34655; // 215
        'h0d8: dout <= -'sd46547; // 216
        'h0d9: dout <=  'sd25865; // 217
        'h0da: dout <=  'sd698; // 218
        'h0db: dout <=  'sd18338; // 219
        'h0dc: dout <= -'sd11444; // 220
        'h0dd: dout <= -'sd25733; // 221
        'h0de: dout <= -'sd17609; // 222
        'h0df: dout <=  'sd56690; // 223
        'h0e0: dout <=  'sd20337; // 224
        'h0e1: dout <=  'sd3077; // 225
        'h0e2: dout <=  'sd7825; // 226
        'h0e3: dout <=  'sd7857; // 227
        'h0e4: dout <=  'sd16888; // 228
        'h0e5: dout <=  'sd48830; // 229
        'h0e6: dout <= -'sd52358; // 230
        'h0e7: dout <=  'sd41092; // 231
        'h0e8: dout <=  'sd8728; // 232
        'h0e9: dout <= -'sd28138; // 233
        'h0ea: dout <= -'sd29361; // 234
        'h0eb: dout <=  'sd27958; // 235
        'h0ec: dout <=  'sd44947; // 236
        'h0ed: dout <=  'sd33131; // 237
        'h0ee: dout <= -'sd45521; // 238
        'h0ef: dout <= -'sd18131; // 239
        'h0f0: dout <=  'sd27013; // 240
        'h0f1: dout <=  'sd30791; // 241
        'h0f2: dout <= -'sd6211; // 242
        'h0f3: dout <=  'sd42643; // 243
        'h0f4: dout <=  'sd35819; // 244
        'h0f5: dout <=  'sd31550; // 245
        'h0f6: dout <=  'sd35691; // 246
        'h0f7: dout <= -'sd21; // 247
        'h0f8: dout <=  'sd44866; // 248
        'h0f9: dout <= -'sd47944; // 249
        'h0fa: dout <=  'sd6034; // 250
        'h0fb: dout <=  'sd21151; // 251
        'h0fc: dout <=  'sd3740; // 252
        'h0fd: dout <=  'sd40435; // 253
        'h0fe: dout <= -'sd48154; // 254
        'h0ff: dout <= -'sd30882; // 255
        'h100: dout <=  'sd16382; // 256
        'h101: dout <=  'sd38167; // 257
        'h102: dout <= -'sd21932; // 258
        'h103: dout <=  'sd24352; // 259
        'h104: dout <= -'sd40899; // 260
        'h105: dout <= -'sd3267; // 261
        'h106: dout <=  'sd49823; // 262
        'h107: dout <= -'sd23102; // 263
        'h108: dout <=  'sd14358; // 264
        'h109: dout <= -'sd48244; // 265
        'h10a: dout <= -'sd56070; // 266
        'h10b: dout <=  'sd16668; // 267
        'h10c: dout <= -'sd25339; // 268
        'h10d: dout <= -'sd25050; // 269
        'h10e: dout <= -'sd5298; // 270
        'h10f: dout <=  'sd14439; // 271
        'h110: dout <=  'sd17103; // 272
        'h111: dout <=  'sd48759; // 273
        'h112: dout <= -'sd42862; // 274
        'h113: dout <=  'sd52244; // 275
        'h114: dout <= -'sd51544; // 276
        'h115: dout <=  'sd41437; // 277
        'h116: dout <=  'sd37893; // 278
        'h117: dout <= -'sd1642; // 279
        'h118: dout <= -'sd21425; // 280
        'h119: dout <= -'sd19344; // 281
        'h11a: dout <= -'sd42584; // 282
        'h11b: dout <= -'sd35506; // 283
        'h11c: dout <= -'sd22355; // 284
        'h11d: dout <=  'sd53286; // 285
        'h11e: dout <=  'sd8849; // 286
        'h11f: dout <= -'sd4281; // 287
        'h120: dout <=  'sd6895; // 288
        'h121: dout <= -'sd13099; // 289
        'h122: dout <= -'sd22818; // 290
        'h123: dout <= -'sd21719; // 291
        'h124: dout <= -'sd6913; // 292
        'h125: dout <=  'sd5049; // 293
        'h126: dout <=  'sd6304; // 294
        'h127: dout <=  'sd31684; // 295
        'h128: dout <= -'sd41590; // 296
        'h129: dout <=  'sd33619; // 297
        'h12a: dout <=  'sd25135; // 298
        'h12b: dout <=  'sd2698; // 299
        'h12c: dout <=  'sd34381; // 300
        'h12d: dout <= -'sd7861; // 301
        'h12e: dout <=  'sd50354; // 302
        'h12f: dout <=  'sd19506; // 303
        'h130: dout <= -'sd44076; // 304
        'h131: dout <= -'sd41947; // 305
        'h132: dout <= -'sd27600; // 306
        'h133: dout <=  'sd35160; // 307
        'h134: dout <=  'sd9875; // 308
        'h135: dout <= -'sd21451; // 309
        'h136: dout <= -'sd2136; // 310
        'h137: dout <= -'sd56322; // 311
        'h138: dout <=  'sd48448; // 312
        'h139: dout <= -'sd33661; // 313
        'h13a: dout <= -'sd38398; // 314
        'h13b: dout <= -'sd38324; // 315
        'h13c: dout <= -'sd33337; // 316
        'h13d: dout <=  'sd20309; // 317
        'h13e: dout <= -'sd18108; // 318
        'h13f: dout <=  'sd21535; // 319
        'h140: dout <=  'sd45289; // 320
        'h141: dout <=  'sd37742; // 321
        'h142: dout <=  'sd17301; // 322
        'h143: dout <= -'sd6692; // 323
        'h144: dout <= -'sd34644; // 324
        'h145: dout <= -'sd15403; // 325
        'h146: dout <= -'sd50383; // 326
        'h147: dout <= -'sd47747; // 327
        'h148: dout <= -'sd38283; // 328
        'h149: dout <=  'sd41325; // 329
        'h14a: dout <=  'sd55549; // 330
        'h14b: dout <=  'sd27784; // 331
        'h14c: dout <= -'sd14853; // 332
        'h14d: dout <= -'sd46922; // 333
        'h14e: dout <=  'sd2853; // 334
        'h14f: dout <=  'sd53018; // 335
        'h150: dout <=  'sd17522; // 336
        'h151: dout <=  'sd13117; // 337
        'h152: dout <= -'sd51437; // 338
        'h153: dout <= -'sd43925; // 339
        'h154: dout <= -'sd40803; // 340
        'h155: dout <= -'sd10919; // 341
        'h156: dout <= -'sd27333; // 342
        'h157: dout <= -'sd29329; // 343
        'h158: dout <= -'sd49274; // 344
        'h159: dout <= -'sd36505; // 345
        'h15a: dout <=  'sd1422; // 346
        'h15b: dout <=  'sd30289; // 347
        'h15c: dout <=  'sd26567; // 348
        'h15d: dout <=  'sd30776; // 349
        'h15e: dout <=  'sd55849; // 350
        'h15f: dout <= -'sd12712; // 351
        'h160: dout <= -'sd36421; // 352
        'h161: dout <=  'sd5274; // 353
        'h162: dout <=  'sd1208; // 354
        'h163: dout <= -'sd51353; // 355
        'h164: dout <= -'sd51367; // 356
        'h165: dout <= -'sd19886; // 357
        'h166: dout <= -'sd56367; // 358
        'h167: dout <=  'sd17202; // 359
        'h168: dout <=  'sd18317; // 360
        'h169: dout <= -'sd12405; // 361
        'h16a: dout <=  'sd48932; // 362
        'h16b: dout <=  'sd20845; // 363
        'h16c: dout <=  'sd17067; // 364
        'h16d: dout <=  'sd26777; // 365
        'h16e: dout <=  'sd31049; // 366
        'h16f: dout <= -'sd9190; // 367
        'h170: dout <= -'sd22816; // 368
        'h171: dout <= -'sd57079; // 369
        'h172: dout <=  'sd4635; // 370
        'h173: dout <=  'sd27807; // 371
        'h174: dout <=  'sd36293; // 372
        'h175: dout <= -'sd6134; // 373
        'h176: dout <=  'sd21722; // 374
        'h177: dout <=  'sd9264; // 375
        'h178: dout <=  'sd29673; // 376
        'h179: dout <=  'sd6547; // 377
        'h17a: dout <=  'sd45297; // 378
        'h17b: dout <=  'sd12851; // 379
        'h17c: dout <= -'sd45062; // 380
        'h17d: dout <=  'sd1358; // 381
        'h17e: dout <=  'sd38706; // 382
        'h17f: dout <= -'sd21351; // 383
        'h180: dout <= -'sd10574; // 384
        'h181: dout <= -'sd45751; // 385
        'h182: dout <= -'sd43264; // 386
        'h183: dout <=  'sd41088; // 387
        'h184: dout <= -'sd20168; // 388
        'h185: dout <=  'sd17170; // 389
        'h186: dout <= -'sd35310; // 390
        'h187: dout <= -'sd15753; // 391
        'h188: dout <= -'sd34425; // 392
        'h189: dout <= -'sd4167; // 393
        'h18a: dout <= -'sd37492; // 394
        'h18b: dout <=  'sd9227; // 395
        'h18c: dout <=  'sd37257; // 396
        'h18d: dout <=  'sd2926; // 397
        'h18e: dout <= -'sd45653; // 398
        'h18f: dout <= -'sd41365; // 399
        'h190: dout <= -'sd3571; // 400
        'h191: dout <= -'sd14122; // 401
        'h192: dout <= -'sd18524; // 402
        'h193: dout <=  'sd56088; // 403
        'h194: dout <= -'sd23803; // 404
        'h195: dout <=  'sd33904; // 405
        'h196: dout <= -'sd22638; // 406
        'h197: dout <= -'sd30832; // 407
        'h198: dout <= -'sd34786; // 408
        'h199: dout <= -'sd49078; // 409
        'h19a: dout <= -'sd33140; // 410
        'h19b: dout <=  'sd22589; // 411
        'h19c: dout <= -'sd5416; // 412
        'h19d: dout <=  'sd28940; // 413
        'h19e: dout <= -'sd54494; // 414
        'h19f: dout <=  'sd27760; // 415
        'h1a0: dout <=  'sd380; // 416
        'h1a1: dout <=  'sd35203; // 417
        'h1a2: dout <= -'sd42462; // 418
        'h1a3: dout <= -'sd27788; // 419
        'h1a4: dout <= -'sd10030; // 420
        'h1a5: dout <= -'sd18007; // 421
        'h1a6: dout <= -'sd45529; // 422
        'h1a7: dout <=  'sd3207; // 423
        'h1a8: dout <=  'sd24132; // 424
        'h1a9: dout <= -'sd51834; // 425
        'h1aa: dout <=  'sd30427; // 426
        'h1ab: dout <=  'sd36488; // 427
        'h1ac: dout <=  'sd48518; // 428
        'h1ad: dout <= -'sd35850; // 429
        'h1ae: dout <= -'sd34333; // 430
        'h1af: dout <=  'sd41894; // 431
        'h1b0: dout <=  'sd9416; // 432
        'h1b1: dout <=  'sd36375; // 433
        'h1b2: dout <=  'sd20015; // 434
        'h1b3: dout <= -'sd49816; // 435
        'h1b4: dout <= -'sd33198; // 436
        'h1b5: dout <=  'sd57084; // 437
        'h1b6: dout <= -'sd47327; // 438
        'h1b7: dout <=  'sd16035; // 439
        'h1b8: dout <=  'sd48699; // 440
        'h1b9: dout <= -'sd19140; // 441
        'h1ba: dout <= -'sd27652; // 442
        'h1bb: dout <=  'sd28232; // 443
        'h1bc: dout <=  'sd15259; // 444
        'h1bd: dout <= -'sd33239; // 445
        'h1be: dout <= -'sd46552; // 446
        'h1bf: dout <= -'sd50696; // 447
        'h1c0: dout <= -'sd32399; // 448
        'h1c1: dout <=  'sd21692; // 449
        'h1c2: dout <=  'sd21456; // 450
        'h1c3: dout <=  'sd35033; // 451
        'h1c4: dout <= -'sd35268; // 452
        'h1c5: dout <= -'sd25828; // 453
        'h1c6: dout <=  'sd8098; // 454
        'h1c7: dout <= -'sd1989; // 455
        'h1c8: dout <=  'sd40963; // 456
        'h1c9: dout <= -'sd44574; // 457
        'h1ca: dout <=  'sd46291; // 458
        'h1cb: dout <= -'sd3227; // 459
        'h1cc: dout <= -'sd24105; // 460
        'h1cd: dout <=  'sd43687; // 461
        'h1ce: dout <= -'sd37472; // 462
        'h1cf: dout <= -'sd24291; // 463
        'h1d0: dout <=  'sd54719; // 464
        'h1d1: dout <=  'sd55105; // 465
        'h1d2: dout <=  'sd1428; // 466
        'h1d3: dout <=  'sd17503; // 467
        'h1d4: dout <=  'sd34594; // 468
        'h1d5: dout <= -'sd13493; // 469
        'h1d6: dout <=  'sd10738; // 470
        'h1d7: dout <= -'sd8923; // 471
        'h1d8: dout <= -'sd35740; // 472
        'h1d9: dout <= -'sd6845; // 473
        'h1da: dout <= -'sd24715; // 474
        'h1db: dout <=  'sd17945; // 475
        'h1dc: dout <= -'sd31327; // 476
        'h1dd: dout <= -'sd10681; // 477
        'h1de: dout <= -'sd54398; // 478
        'h1df: dout <= -'sd44092; // 479
        'h1e0: dout <=  'sd24361; // 480
        'h1e1: dout <= -'sd41903; // 481
        'h1e2: dout <= -'sd49749; // 482
        'h1e3: dout <= -'sd45126; // 483
        'h1e4: dout <=  'sd26449; // 484
        'h1e5: dout <= -'sd26921; // 485
        'h1e6: dout <=  'sd29139; // 486
        'h1e7: dout <= -'sd25958; // 487
        'h1e8: dout <= -'sd11716; // 488
        'h1e9: dout <= -'sd40696; // 489
        'h1ea: dout <= -'sd25152; // 490
        'h1eb: dout <=  'sd18891; // 491
        'h1ec: dout <= -'sd1765; // 492
        'h1ed: dout <= -'sd28121; // 493
        'h1ee: dout <=  'sd47592; // 494
        'h1ef: dout <=  'sd49414; // 495
        'h1f0: dout <=  'sd38314; // 496
        'h1f1: dout <= -'sd1019; // 497
        'h1f2: dout <= -'sd2506; // 498
        'h1f3: dout <=  'sd16694; // 499
        'h1f4: dout <= -'sd54505; // 500
        'h1f5: dout <=  'sd21101; // 501
        'h1f6: dout <= -'sd54732; // 502
        'h1f7: dout <= -'sd30954; // 503
        'h1f8: dout <= -'sd20164; // 504
        'h1f9: dout <=  'sd32431; // 505
        'h1fa: dout <= -'sd6234; // 506
        'h1fb: dout <=  'sd34659; // 507
        'h1fc: dout <= -'sd25543; // 508
        'h1fd: dout <= -'sd42928; // 509
        'h1fe: dout <=  'sd3226; // 510
        'h1ff: dout <= -'sd43959; // 511
        'h200: dout <=  'sd14026; // 512
        'h201: dout <=  'sd56152; // 513
        'h202: dout <=  'sd19056; // 514
        'h203: dout <= -'sd47498; // 515
        'h204: dout <= -'sd10420; // 516
        'h205: dout <= -'sd20446; // 517
        'h206: dout <=  'sd1155; // 518
        'h207: dout <=  'sd8793; // 519
        'h208: dout <=  'sd11564; // 520
        'h209: dout <=  'sd41291; // 521
        'h20a: dout <=  'sd50333; // 522
        'h20b: dout <= -'sd55309; // 523
        'h20c: dout <=  'sd8264; // 524
        'h20d: dout <= -'sd14291; // 525
        'h20e: dout <= -'sd26159; // 526
        'h20f: dout <= -'sd14825; // 527
        'h210: dout <= -'sd49709; // 528
        'h211: dout <= -'sd20012; // 529
        'h212: dout <= -'sd49838; // 530
        'h213: dout <=  'sd5962; // 531
        'h214: dout <=  'sd12755; // 532
        'h215: dout <=  'sd23303; // 533
        'h216: dout <=  'sd21303; // 534
        'h217: dout <=  'sd9211; // 535
        'h218: dout <= -'sd54628; // 536
        'h219: dout <=  'sd6216; // 537
        'h21a: dout <= -'sd34724; // 538
        'h21b: dout <=  'sd36950; // 539
        'h21c: dout <= -'sd37049; // 540
        'h21d: dout <= -'sd16934; // 541
        'h21e: dout <=  'sd8698; // 542
        'h21f: dout <= -'sd48489; // 543
        'h220: dout <=  'sd7171; // 544
        'h221: dout <=  'sd23174; // 545
        'h222: dout <= -'sd12859; // 546
        'h223: dout <= -'sd2239; // 547
        'h224: dout <= -'sd31227; // 548
        'h225: dout <= -'sd51068; // 549
        'h226: dout <= -'sd40023; // 550
        'h227: dout <= -'sd52055; // 551
        'h228: dout <=  'sd1760; // 552
        'h229: dout <= -'sd23532; // 553
        'h22a: dout <=  'sd43312; // 554
        'h22b: dout <=  'sd50134; // 555
        'h22c: dout <=  'sd38023; // 556
        'h22d: dout <= -'sd32169; // 557
        'h22e: dout <= -'sd21917; // 558
        'h22f: dout <= -'sd16207; // 559
        'h230: dout <= -'sd11205; // 560
        'h231: dout <= -'sd10931; // 561
        'h232: dout <= -'sd13850; // 562
        'h233: dout <= -'sd17530; // 563
        'h234: dout <= -'sd14942; // 564
        'h235: dout <= -'sd52960; // 565
        'h236: dout <=  'sd12130; // 566
        'h237: dout <=  'sd36644; // 567
        'h238: dout <= -'sd9607; // 568
        'h239: dout <= -'sd39615; // 569
        'h23a: dout <=  'sd12984; // 570
        'h23b: dout <=  'sd32104; // 571
        'h23c: dout <= -'sd45565; // 572
        'h23d: dout <= -'sd31759; // 573
        'h23e: dout <= -'sd40713; // 574
        'h23f: dout <=  'sd52508; // 575
        'h240: dout <=  'sd39277; // 576
        'h241: dout <= -'sd18944; // 577
        'h242: dout <= -'sd14688; // 578
        'h243: dout <= -'sd20164; // 579
        'h244: dout <=  'sd37518; // 580
        'h245: dout <= -'sd42848; // 581
        'h246: dout <=  'sd12645; // 582
        'h247: dout <=  'sd28120; // 583
        'h248: dout <=  'sd35930; // 584
        'h249: dout <=  'sd9669; // 585
        'h24a: dout <= -'sd42954; // 586
        'h24b: dout <= -'sd10479; // 587
        'h24c: dout <= -'sd31323; // 588
        'h24d: dout <= -'sd10947; // 589
        'h24e: dout <= -'sd33375; // 590
        'h24f: dout <= -'sd26264; // 591
        'h250: dout <= -'sd51191; // 592
        'h251: dout <=  'sd36289; // 593
        'h252: dout <= -'sd35968; // 594
        'h253: dout <=  'sd45463; // 595
        'h254: dout <=  'sd9764; // 596
        'h255: dout <=  'sd20771; // 597
        'h256: dout <= -'sd21980; // 598
        'h257: dout <= -'sd53503; // 599
        'h258: dout <= -'sd9669; // 600
        'h259: dout <=  'sd43505; // 601
        'h25a: dout <= -'sd37532; // 602
        'h25b: dout <= -'sd46934; // 603
        'h25c: dout <= -'sd41784; // 604
        'h25d: dout <=  'sd5750; // 605
        'h25e: dout <= -'sd529; // 606
        'h25f: dout <= -'sd18425; // 607
        'h260: dout <=  'sd1586; // 608
        'h261: dout <= -'sd46369; // 609
        'h262: dout <= -'sd7428; // 610
        'h263: dout <= -'sd14980; // 611
        'h264: dout <=  'sd16287; // 612
        'h265: dout <=  'sd4432; // 613
        'h266: dout <=  'sd4096; // 614
        'h267: dout <= -'sd25760; // 615
        'h268: dout <= -'sd11455; // 616
        'h269: dout <=  'sd41883; // 617
        'h26a: dout <= -'sd20045; // 618
        'h26b: dout <= -'sd13637; // 619
        'h26c: dout <=  'sd29009; // 620
        'h26d: dout <=  'sd42981; // 621
        'h26e: dout <=  'sd23738; // 622
        'h26f: dout <= -'sd57083; // 623
        'h270: dout <=  'sd42448; // 624
        'h271: dout <= -'sd48972; // 625
        'h272: dout <= -'sd42822; // 626
        'h273: dout <= -'sd49932; // 627
        'h274: dout <=  'sd1455; // 628
        'h275: dout <= -'sd28327; // 629
        'h276: dout <= -'sd3346; // 630
        'h277: dout <= -'sd27416; // 631
        'h278: dout <= -'sd54758; // 632
        'h279: dout <=  'sd2443; // 633
        'h27a: dout <= -'sd22812; // 634
        'h27b: dout <= -'sd27585; // 635
        'h27c: dout <=  'sd2555; // 636
        'h27d: dout <= -'sd619; // 637
        'h27e: dout <=  'sd56755; // 638
        'h27f: dout <=  'sd25159; // 639
        'h280: dout <=  'sd48938; // 640
        'h281: dout <=  'sd4601; // 641
        'h282: dout <=  'sd43343; // 642
        'h283: dout <=  'sd53876; // 643
        'h284: dout <= -'sd49349; // 644
        'h285: dout <=  'sd38669; // 645
        'h286: dout <=  'sd56051; // 646
        'h287: dout <= -'sd17913; // 647
        'h288: dout <= -'sd9935; // 648
        'h289: dout <=  'sd51989; // 649
        'h28a: dout <= -'sd3450; // 650
        'h28b: dout <=  'sd46683; // 651
        'h28c: dout <= -'sd5896; // 652
        'h28d: dout <= -'sd19084; // 653
        'h28e: dout <=  'sd38134; // 654
        'h28f: dout <= -'sd6327; // 655
        'h290: dout <= -'sd42169; // 656
        'h291: dout <= -'sd26323; // 657
        'h292: dout <= -'sd50115; // 658
        'h293: dout <= -'sd51218; // 659
        'h294: dout <= -'sd43605; // 660
        'h295: dout <=  'sd10715; // 661
        'h296: dout <= -'sd36658; // 662
        'h297: dout <= -'sd14205; // 663
        'h298: dout <= -'sd23555; // 664
        'h299: dout <=  'sd16577; // 665
        'h29a: dout <= -'sd12871; // 666
        'h29b: dout <=  'sd57093; // 667
        'h29c: dout <=  'sd41193; // 668
        'h29d: dout <=  'sd31688; // 669
        'h29e: dout <= -'sd52924; // 670
        'h29f: dout <= -'sd52650; // 671
        'h2a0: dout <= -'sd49388; // 672
        'h2a1: dout <= -'sd500; // 673
        'h2a2: dout <= -'sd18188; // 674
        'h2a3: dout <=  'sd29286; // 675
        'h2a4: dout <= -'sd30110; // 676
        'h2a5: dout <= -'sd11978; // 677
        'h2a6: dout <= -'sd1643; // 678
        'h2a7: dout <=  'sd5475; // 679
        'h2a8: dout <=  'sd51761; // 680
        'h2a9: dout <= -'sd35441; // 681
        'h2aa: dout <= -'sd1820; // 682
        'h2ab: dout <= -'sd2648; // 683
        'h2ac: dout <=  'sd25091; // 684
        'h2ad: dout <= -'sd25532; // 685
        'h2ae: dout <=  'sd22481; // 686
        'h2af: dout <=  'sd24309; // 687
        'h2b0: dout <=  'sd18213; // 688
        'h2b1: dout <=  'sd49902; // 689
        'h2b2: dout <= -'sd9886; // 690
        'h2b3: dout <= -'sd50846; // 691
        'h2b4: dout <=  'sd11432; // 692
        'h2b5: dout <=  'sd5117; // 693
        'h2b6: dout <=  'sd18885; // 694
        'h2b7: dout <= -'sd1634; // 695
        'h2b8: dout <=  'sd574; // 696
        'h2b9: dout <=  'sd40438; // 697
        'h2ba: dout <= -'sd4724; // 698
        'h2bb: dout <=  'sd39209; // 699
        'h2bc: dout <=  'sd33887; // 700
        'h2bd: dout <= -'sd52896; // 701
        'h2be: dout <=  'sd33108; // 702
        'h2bf: dout <= -'sd9467; // 703
        'h2c0: dout <= -'sd47003; // 704
        'h2c1: dout <= -'sd35904; // 705
        'h2c2: dout <=  'sd40353; // 706
        'h2c3: dout <=  'sd16715; // 707
        'h2c4: dout <=  'sd6217; // 708
        'h2c5: dout <=  'sd897; // 709
        'h2c6: dout <= -'sd45686; // 710
        'h2c7: dout <=  'sd23570; // 711
        'h2c8: dout <= -'sd4434; // 712
        'h2c9: dout <= -'sd43489; // 713
        'h2ca: dout <=  'sd9849; // 714
        'h2cb: dout <= -'sd25966; // 715
        'h2cc: dout <=  'sd50146; // 716
        'h2cd: dout <= -'sd16867; // 717
        'h2ce: dout <=  'sd34760; // 718
        'h2cf: dout <=  'sd45842; // 719
        'h2d0: dout <= -'sd38683; // 720
        'h2d1: dout <=  'sd27880; // 721
        'h2d2: dout <= -'sd38655; // 722
        'h2d3: dout <= -'sd42119; // 723
        'h2d4: dout <= -'sd34266; // 724
        'h2d5: dout <=  'sd21285; // 725
        'h2d6: dout <= -'sd40518; // 726
        'h2d7: dout <=  'sd39808; // 727
        'h2d8: dout <= -'sd49961; // 728
        'h2d9: dout <= -'sd16854; // 729
        'h2da: dout <=  'sd40554; // 730
        'h2db: dout <= -'sd23852; // 731
        'h2dc: dout <=  'sd54970; // 732
        'h2dd: dout <=  'sd25373; // 733
        'h2de: dout <=  'sd20866; // 734
        'h2df: dout <=  'sd21056; // 735
        'h2e0: dout <=  'sd34082; // 736
        'h2e1: dout <=  'sd13272; // 737
        'h2e2: dout <= -'sd48060; // 738
        'h2e3: dout <= -'sd26970; // 739
        'h2e4: dout <=  'sd22128; // 740
        'h2e5: dout <= -'sd24720; // 741
        'h2e6: dout <=  'sd54376; // 742
        'h2e7: dout <=  'sd35182; // 743
        'h2e8: dout <=  'sd14747; // 744
        'h2e9: dout <= -'sd41723; // 745
        'h2ea: dout <=  'sd51783; // 746
        'h2eb: dout <= -'sd10927; // 747
        'h2ec: dout <=  'sd28394; // 748
        'h2ed: dout <= -'sd22; // 749
        'h2ee: dout <=  'sd49363; // 750
        'h2ef: dout <= -'sd50243; // 751
        'h2f0: dout <= -'sd35032; // 752
        'h2f1: dout <= -'sd50942; // 753
        'h2f2: dout <= -'sd3751; // 754
        'h2f3: dout <= -'sd15784; // 755
        'h2f4: dout <=  'sd33041; // 756
        'h2f5: dout <=  'sd18878; // 757
        'h2f6: dout <=  'sd55873; // 758
        'h2f7: dout <=  'sd20527; // 759
        'h2f8: dout <=  'sd39258; // 760
        'h2f9: dout <= -'sd51541; // 761
        'h2fa: dout <= -'sd16124; // 762
        'h2fb: dout <=  'sd12867; // 763
        'h2fc: dout <=  'sd15275; // 764
        'h2fd: dout <=  'sd41938; // 765
        'h2fe: dout <= -'sd13032; // 766
        'h2ff: dout <=  'sd11455; // 767
        'h300: dout <= -'sd41919; // 768
        'h301: dout <=  'sd47313; // 769
        'h302: dout <=  'sd43295; // 770
        'h303: dout <= -'sd30037; // 771
        'h304: dout <=  'sd5237; // 772
        'h305: dout <=  'sd45912; // 773
        'h306: dout <= -'sd37990; // 774
        'h307: dout <= -'sd56670; // 775
        'h308: dout <=  'sd55076; // 776
        'h309: dout <=  'sd29124; // 777
        'h30a: dout <= -'sd42368; // 778
        'h30b: dout <= -'sd54574; // 779
        'h30c: dout <=  'sd9057; // 780
        'h30d: dout <=  'sd49299; // 781
        'h30e: dout <= -'sd30298; // 782
        'h30f: dout <= -'sd8257; // 783
        'h310: dout <= -'sd43704; // 784
        'h311: dout <=  'sd22814; // 785
        'h312: dout <= -'sd2353; // 786
        'h313: dout <=  'sd43001; // 787
        'h314: dout <=  'sd5244; // 788
        'h315: dout <= -'sd13250; // 789
        'h316: dout <=  'sd15465; // 790
        'h317: dout <= -'sd30598; // 791
        'h318: dout <=  'sd29829; // 792
        'h319: dout <=  'sd56742; // 793
        'h31a: dout <= -'sd57026; // 794
        'h31b: dout <=  'sd41038; // 795
        'h31c: dout <=  'sd21324; // 796
        'h31d: dout <=  'sd13928; // 797
        'h31e: dout <=  'sd42770; // 798
        'h31f: dout <=  'sd43745; // 799
        'h320: dout <=  'sd48583; // 800
        'h321: dout <=  'sd36116; // 801
        'h322: dout <= -'sd23591; // 802
        'h323: dout <=  'sd33401; // 803
        'h324: dout <=  'sd28422; // 804
        'h325: dout <=  'sd46511; // 805
        'h326: dout <= -'sd54645; // 806
        'h327: dout <=  'sd48035; // 807
        'h328: dout <=  'sd6878; // 808
        'h329: dout <= -'sd14004; // 809
        'h32a: dout <= -'sd4869; // 810
        'h32b: dout <= -'sd1649; // 811
        'h32c: dout <=  'sd43622; // 812
        'h32d: dout <=  'sd44569; // 813
        'h32e: dout <= -'sd7097; // 814
        'h32f: dout <= -'sd34222; // 815
        'h330: dout <=  'sd24122; // 816
        'h331: dout <= -'sd54570; // 817
        'h332: dout <=  'sd2347; // 818
        'h333: dout <= -'sd45226; // 819
        'h334: dout <=  'sd44841; // 820
        'h335: dout <= -'sd15559; // 821
        'h336: dout <= -'sd44616; // 822
        'h337: dout <=  'sd47650; // 823
        'h338: dout <=  'sd27671; // 824
        'h339: dout <=  'sd48884; // 825
        'h33a: dout <= -'sd31346; // 826
        'h33b: dout <= -'sd28505; // 827
        'h33c: dout <=  'sd34313; // 828
        'h33d: dout <= -'sd27849; // 829
        'h33e: dout <=  'sd11138; // 830
        'h33f: dout <= -'sd4304; // 831
        'h340: dout <= -'sd41462; // 832
        'h341: dout <= -'sd6365; // 833
        'h342: dout <= -'sd47569; // 834
        'h343: dout <=  'sd45497; // 835
        'h344: dout <=  'sd44049; // 836
        'h345: dout <= -'sd6677; // 837
        'h346: dout <= -'sd36303; // 838
        'h347: dout <= -'sd17145; // 839
        'h348: dout <=  'sd40068; // 840
        'h349: dout <= -'sd14180; // 841
        'h34a: dout <= -'sd182; // 842
        'h34b: dout <= -'sd18797; // 843
        'h34c: dout <= -'sd37252; // 844
        'h34d: dout <= -'sd56226; // 845
        'h34e: dout <= -'sd29568; // 846
        'h34f: dout <=  'sd36354; // 847
        'h350: dout <= -'sd42735; // 848
        'h351: dout <= -'sd49074; // 849
        'h352: dout <=  'sd17572; // 850
        'h353: dout <=  'sd38162; // 851
        'h354: dout <=  'sd36843; // 852
        'h355: dout <= -'sd24136; // 853
        'h356: dout <=  'sd55049; // 854
        'h357: dout <=  'sd15356; // 855
        'h358: dout <=  'sd48368; // 856
        'h359: dout <=  'sd44757; // 857
        'h35a: dout <=  'sd1590; // 858
        'h35b: dout <= -'sd51286; // 859
        'h35c: dout <= -'sd13033; // 860
        'h35d: dout <= -'sd12950; // 861
        'h35e: dout <=  'sd49573; // 862
        'h35f: dout <= -'sd23517; // 863
        'h360: dout <= -'sd48820; // 864
        'h361: dout <=  'sd6099; // 865
        'h362: dout <=  'sd24982; // 866
        'h363: dout <= -'sd63; // 867
        'h364: dout <=  'sd52705; // 868
        'h365: dout <= -'sd47573; // 869
        'h366: dout <= -'sd54127; // 870
        'h367: dout <=  'sd30408; // 871
        'h368: dout <=  'sd22230; // 872
        'h369: dout <=  'sd8258; // 873
        'h36a: dout <=  'sd46725; // 874
        'h36b: dout <=  'sd51548; // 875
        'h36c: dout <=  'sd19687; // 876
        'h36d: dout <=  'sd10939; // 877
        'h36e: dout <=  'sd21009; // 878
        'h36f: dout <= -'sd32776; // 879
        'h370: dout <=  'sd4672; // 880
        'h371: dout <=  'sd7573; // 881
        'h372: dout <= -'sd15245; // 882
        'h373: dout <=  'sd3884; // 883
        'h374: dout <=  'sd26240; // 884
        'h375: dout <=  'sd56735; // 885
        'h376: dout <=  'sd47685; // 886
        'h377: dout <= -'sd11468; // 887
        'h378: dout <=  'sd2609; // 888
        'h379: dout <= -'sd33858; // 889
        'h37a: dout <=  'sd29307; // 890
        'h37b: dout <=  'sd48743; // 891
        'h37c: dout <=  'sd48438; // 892
        'h37d: dout <= -'sd51137; // 893
        'h37e: dout <= -'sd787; // 894
        'h37f: dout <=  'sd5683; // 895
        'h380: dout <= -'sd43247; // 896
        'h381: dout <=  'sd22832; // 897
        'h382: dout <=  'sd6573; // 898
        'h383: dout <=  'sd36173; // 899
        'h384: dout <=  'sd26464; // 900
        'h385: dout <=  'sd21060; // 901
        'h386: dout <=  'sd20846; // 902
        'h387: dout <= -'sd20793; // 903
        'h388: dout <= -'sd22452; // 904
        'h389: dout <= -'sd54740; // 905
        'h38a: dout <=  'sd10749; // 906
        'h38b: dout <=  'sd12956; // 907
        'h38c: dout <= -'sd35739; // 908
        'h38d: dout <= -'sd11468; // 909
        'h38e: dout <=  'sd26176; // 910
        'h38f: dout <=  'sd50283; // 911
        'h390: dout <= -'sd12197; // 912
        'h391: dout <= -'sd6584; // 913
        'h392: dout <=  'sd50021; // 914
        'h393: dout <= -'sd23374; // 915
        'h394: dout <= -'sd45425; // 916
        'h395: dout <= -'sd1746; // 917
        'h396: dout <=  'sd35997; // 918
        'h397: dout <=  'sd25416; // 919
        'h398: dout <=  'sd39104; // 920
        'h399: dout <= -'sd40312; // 921
        'h39a: dout <= -'sd17216; // 922
        'h39b: dout <=  'sd38190; // 923
        'h39c: dout <=  'sd34863; // 924
        'h39d: dout <=  'sd53986; // 925
        'h39e: dout <= -'sd38286; // 926
        'h39f: dout <=  'sd7839; // 927
        'h3a0: dout <= -'sd37388; // 928
        'h3a1: dout <= -'sd7053; // 929
        'h3a2: dout <=  'sd39347; // 930
        'h3a3: dout <=  'sd52194; // 931
        'h3a4: dout <=  'sd20237; // 932
        'h3a5: dout <= -'sd25310; // 933
        'h3a6: dout <=  'sd12061; // 934
        'h3a7: dout <= -'sd30802; // 935
        'h3a8: dout <= -'sd55402; // 936
        'h3a9: dout <= -'sd28781; // 937
        'h3aa: dout <= -'sd35813; // 938
        'h3ab: dout <= -'sd28021; // 939
        'h3ac: dout <= -'sd16943; // 940
        'h3ad: dout <=  'sd3715; // 941
        'h3ae: dout <=  'sd22134; // 942
        'h3af: dout <=  'sd1127; // 943
        'h3b0: dout <=  'sd15901; // 944
        'h3b1: dout <= -'sd35039; // 945
        'h3b2: dout <= -'sd22638; // 946
        'h3b3: dout <= -'sd16025; // 947
        'h3b4: dout <=  'sd31679; // 948
        'h3b5: dout <= -'sd53604; // 949
        'h3b6: dout <= -'sd4214; // 950
        'h3b7: dout <= -'sd8794; // 951
        'h3b8: dout <=  'sd32649; // 952
        'h3b9: dout <=  'sd47639; // 953
        'h3ba: dout <= -'sd50459; // 954
        'h3bb: dout <= -'sd29516; // 955
        'h3bc: dout <=  'sd2040; // 956
        'h3bd: dout <=  'sd46870; // 957
        'h3be: dout <=  'sd13546; // 958
        'h3bf: dout <= -'sd21204; // 959
        'h3c0: dout <= -'sd45215; // 960
        'h3c1: dout <= -'sd2664; // 961
        'h3c2: dout <= -'sd57086; // 962
        'h3c3: dout <= -'sd10617; // 963
        'h3c4: dout <= -'sd1275; // 964
        'h3c5: dout <= -'sd21471; // 965
        'h3c6: dout <= -'sd40972; // 966
        'h3c7: dout <= -'sd43618; // 967
        'h3c8: dout <=  'sd46732; // 968
        'h3c9: dout <=  'sd20311; // 969
        'h3ca: dout <=  'sd57342; // 970
        'h3cb: dout <=  'sd32373; // 971
        'h3cc: dout <= -'sd18075; // 972
        'h3cd: dout <=  'sd19234; // 973
        'h3ce: dout <= -'sd3989; // 974
        'h3cf: dout <= -'sd45971; // 975
        'h3d0: dout <=  'sd39860; // 976
        'h3d1: dout <= -'sd48197; // 977
        'h3d2: dout <= -'sd7128; // 978
        'h3d3: dout <= -'sd37539; // 979
        'h3d4: dout <=  'sd9933; // 980
        'h3d5: dout <=  'sd33656; // 981
        'h3d6: dout <= -'sd17333; // 982
        'h3d7: dout <=  'sd17679; // 983
        'h3d8: dout <= -'sd53712; // 984
        'h3d9: dout <= -'sd45694; // 985
        'h3da: dout <=  'sd10126; // 986
        'h3db: dout <= -'sd17961; // 987
        'h3dc: dout <= -'sd8978; // 988
        'h3dd: dout <=  'sd46837; // 989
        'h3de: dout <=  'sd6470; // 990
        'h3df: dout <=  'sd23163; // 991
        'h3e0: dout <=  'sd48083; // 992
        'h3e1: dout <= -'sd10829; // 993
        'h3e2: dout <= -'sd18280; // 994
        'h3e3: dout <=  'sd40941; // 995
        'h3e4: dout <= -'sd10202; // 996
        'h3e5: dout <=  'sd17593; // 997
        'h3e6: dout <=  'sd21765; // 998
        'h3e7: dout <=  'sd8224; // 999
        'h3e8: dout <= -'sd24265; // 1000
        'h3e9: dout <= -'sd49719; // 1001
        'h3ea: dout <=  'sd29607; // 1002
        'h3eb: dout <=  'sd13901; // 1003
        'h3ec: dout <= -'sd52986; // 1004
        'h3ed: dout <=  'sd9843; // 1005
        'h3ee: dout <=  'sd27589; // 1006
        'h3ef: dout <=  'sd7609; // 1007
        'h3f0: dout <=  'sd54962; // 1008
        'h3f1: dout <=  'sd17719; // 1009
        'h3f2: dout <= -'sd48559; // 1010
        'h3f3: dout <= -'sd6388; // 1011
        'h3f4: dout <= -'sd52782; // 1012
        'h3f5: dout <=  'sd13435; // 1013
        'h3f6: dout <= -'sd28153; // 1014
        'h3f7: dout <=  'sd44842; // 1015
        'h3f8: dout <= -'sd561; // 1016
        'h3f9: dout <= -'sd15294; // 1017
        'h3fa: dout <= -'sd17213; // 1018
        'h3fb: dout <= -'sd19998; // 1019
        'h3fc: dout <=  'sd24801; // 1020
        'h3fd: dout <=  'sd31980; // 1021
        'h3fe: dout <= -'sd5828; // 1022
        'h3ff: dout <= -'sd38985; // 1023
        'h400: dout <=  'sd43154; // 1024
        'h401: dout <=  'sd53983; // 1025
        'h402: dout <= -'sd25772; // 1026
        'h403: dout <= -'sd46145; // 1027
        'h404: dout <=  'sd38117; // 1028
        'h405: dout <=  'sd3509; // 1029
        'h406: dout <= -'sd43171; // 1030
        'h407: dout <= -'sd16667; // 1031
        'h408: dout <= -'sd7889; // 1032
        'h409: dout <=  'sd46701; // 1033
        'h40a: dout <= -'sd49409; // 1034
        'h40b: dout <=  'sd12109; // 1035
        'h40c: dout <=  'sd41584; // 1036
        'h40d: dout <=  'sd33075; // 1037
        'h40e: dout <=  'sd40468; // 1038
        'h40f: dout <=  'sd52953; // 1039
        'h410: dout <=  'sd33352; // 1040
        'h411: dout <= -'sd38913; // 1041
        'h412: dout <= -'sd42491; // 1042
        'h413: dout <=  'sd8306; // 1043
        'h414: dout <=  'sd3047; // 1044
        'h415: dout <= -'sd54383; // 1045
        'h416: dout <= -'sd24598; // 1046
        'h417: dout <= -'sd41194; // 1047
        'h418: dout <=  'sd2322; // 1048
        'h419: dout <=  'sd25527; // 1049
        'h41a: dout <= -'sd20800; // 1050
        'h41b: dout <=  'sd31884; // 1051
        'h41c: dout <=  'sd30077; // 1052
        'h41d: dout <=  'sd54428; // 1053
        'h41e: dout <=  'sd31100; // 1054
        'h41f: dout <=  'sd16437; // 1055
        'h420: dout <= -'sd20958; // 1056
        'h421: dout <=  'sd17865; // 1057
        'h422: dout <=  'sd20968; // 1058
        'h423: dout <= -'sd33916; // 1059
        'h424: dout <= -'sd48458; // 1060
        'h425: dout <= -'sd31566; // 1061
        'h426: dout <=  'sd14366; // 1062
        'h427: dout <=  'sd12244; // 1063
        'h428: dout <=  'sd43264; // 1064
        'h429: dout <=  'sd29161; // 1065
        'h42a: dout <= -'sd4906; // 1066
        'h42b: dout <= -'sd28483; // 1067
        'h42c: dout <= -'sd51753; // 1068
        'h42d: dout <= -'sd30932; // 1069
        'h42e: dout <=  'sd39744; // 1070
        'h42f: dout <=  'sd54747; // 1071
        'h430: dout <=  'sd37403; // 1072
        'h431: dout <= -'sd40809; // 1073
        'h432: dout <=  'sd32192; // 1074
        'h433: dout <=  'sd29132; // 1075
        'h434: dout <=  'sd10866; // 1076
        'h435: dout <= -'sd7401; // 1077
        'h436: dout <=  'sd27035; // 1078
        'h437: dout <=  'sd5801; // 1079
        'h438: dout <= -'sd11578; // 1080
        'h439: dout <= -'sd3944; // 1081
        'h43a: dout <= -'sd24550; // 1082
        'h43b: dout <=  'sd9162; // 1083
        'h43c: dout <= -'sd42733; // 1084
        'h43d: dout <=  'sd43240; // 1085
        'h43e: dout <=  'sd42968; // 1086
        'h43f: dout <= -'sd1204; // 1087
        'h440: dout <= -'sd13169; // 1088
        'h441: dout <= -'sd41071; // 1089
        'h442: dout <=  'sd9688; // 1090
        'h443: dout <= -'sd2426; // 1091
        'h444: dout <= -'sd55561; // 1092
        'h445: dout <=  'sd56043; // 1093
        'h446: dout <=  'sd53934; // 1094
        'h447: dout <= -'sd47380; // 1095
        'h448: dout <= -'sd42631; // 1096
        'h449: dout <= -'sd43213; // 1097
        'h44a: dout <=  'sd25522; // 1098
        'h44b: dout <=  'sd22265; // 1099
        'h44c: dout <=  'sd2342; // 1100
        'h44d: dout <=  'sd5733; // 1101
        'h44e: dout <= -'sd56025; // 1102
        'h44f: dout <= -'sd28179; // 1103
        'h450: dout <=  'sd38450; // 1104
        'h451: dout <=  'sd17187; // 1105
        'h452: dout <= -'sd10693; // 1106
        'h453: dout <= -'sd32844; // 1107
        'h454: dout <=  'sd49903; // 1108
        'h455: dout <= -'sd15736; // 1109
        'h456: dout <= -'sd9855; // 1110
        'h457: dout <= -'sd36077; // 1111
        'h458: dout <= -'sd5748; // 1112
        'h459: dout <=  'sd42022; // 1113
        'h45a: dout <= -'sd24527; // 1114
        'h45b: dout <= -'sd4673; // 1115
        'h45c: dout <=  'sd20489; // 1116
        'h45d: dout <= -'sd24101; // 1117
        'h45e: dout <=  'sd1547; // 1118
        'h45f: dout <=  'sd5747; // 1119
        'h460: dout <= -'sd22642; // 1120
        'h461: dout <=  'sd6835; // 1121
        'h462: dout <= -'sd13662; // 1122
        'h463: dout <= -'sd16957; // 1123
        'h464: dout <= -'sd8562; // 1124
        'h465: dout <=  'sd14042; // 1125
        'h466: dout <= -'sd4664; // 1126
        'h467: dout <=  'sd33678; // 1127
        'h468: dout <=  'sd41380; // 1128
        'h469: dout <=  'sd55819; // 1129
        'h46a: dout <=  'sd1649; // 1130
        'h46b: dout <=  'sd7093; // 1131
        'h46c: dout <= -'sd9776; // 1132
        'h46d: dout <= -'sd38966; // 1133
        'h46e: dout <= -'sd26760; // 1134
        'h46f: dout <=  'sd52076; // 1135
        'h470: dout <=  'sd17942; // 1136
        'h471: dout <=  'sd26778; // 1137
        'h472: dout <=  'sd55852; // 1138
        'h473: dout <=  'sd12929; // 1139
        'h474: dout <=  'sd54725; // 1140
        'h475: dout <=  'sd1630; // 1141
        'h476: dout <=  'sd34370; // 1142
        'h477: dout <=  'sd11435; // 1143
        'h478: dout <= -'sd8606; // 1144
        'h479: dout <= -'sd7419; // 1145
        'h47a: dout <= -'sd10876; // 1146
        'h47b: dout <= -'sd41839; // 1147
        'h47c: dout <= -'sd7667; // 1148
        'h47d: dout <=  'sd37858; // 1149
        'h47e: dout <= -'sd4591; // 1150
        'h47f: dout <= -'sd14078; // 1151
        'h480: dout <=  'sd21887; // 1152
        'h481: dout <= -'sd25253; // 1153
        'h482: dout <=  'sd8615; // 1154
        'h483: dout <= -'sd21556; // 1155
        'h484: dout <= -'sd53935; // 1156
        'h485: dout <= -'sd43175; // 1157
        'h486: dout <= -'sd13877; // 1158
        'h487: dout <= -'sd53547; // 1159
        'h488: dout <=  'sd21936; // 1160
        'h489: dout <= -'sd21612; // 1161
        'h48a: dout <=  'sd42849; // 1162
        'h48b: dout <=  'sd36210; // 1163
        'h48c: dout <= -'sd28174; // 1164
        'h48d: dout <= -'sd41029; // 1165
        'h48e: dout <=  'sd56977; // 1166
        'h48f: dout <=  'sd13867; // 1167
        'h490: dout <=  'sd8425; // 1168
        'h491: dout <=  'sd56315; // 1169
        'h492: dout <=  'sd456; // 1170
        'h493: dout <= -'sd17566; // 1171
        'h494: dout <=  'sd19151; // 1172
        'h495: dout <= -'sd26407; // 1173
        'h496: dout <= -'sd43889; // 1174
        'h497: dout <=  'sd54233; // 1175
        'h498: dout <= -'sd26551; // 1176
        'h499: dout <=  'sd27988; // 1177
        'h49a: dout <= -'sd45881; // 1178
        'h49b: dout <=  'sd53635; // 1179
        'h49c: dout <= -'sd16827; // 1180
        'h49d: dout <= -'sd14494; // 1181
        'h49e: dout <= -'sd54311; // 1182
        'h49f: dout <= -'sd41435; // 1183
        'h4a0: dout <= -'sd2484; // 1184
        'h4a1: dout <= -'sd51319; // 1185
        'h4a2: dout <= -'sd51836; // 1186
        'h4a3: dout <= -'sd47156; // 1187
        'h4a4: dout <= -'sd45271; // 1188
        'h4a5: dout <= -'sd2421; // 1189
        'h4a6: dout <=  'sd14339; // 1190
        'h4a7: dout <= -'sd20732; // 1191
        'h4a8: dout <=  'sd15839; // 1192
        'h4a9: dout <= -'sd27455; // 1193
        'h4aa: dout <=  'sd25145; // 1194
        'h4ab: dout <= -'sd5382; // 1195
        'h4ac: dout <=  'sd48624; // 1196
        'h4ad: dout <= -'sd31683; // 1197
        'h4ae: dout <= -'sd40735; // 1198
        'h4af: dout <= -'sd20897; // 1199
        'h4b0: dout <=  'sd2688; // 1200
        'h4b1: dout <= -'sd42295; // 1201
        'h4b2: dout <=  'sd9179; // 1202
        'h4b3: dout <=  'sd20501; // 1203
        'h4b4: dout <= -'sd56314; // 1204
        'h4b5: dout <= -'sd13629; // 1205
        'h4b6: dout <=  'sd52192; // 1206
        'h4b7: dout <=  'sd7149; // 1207
        'h4b8: dout <= -'sd26431; // 1208
        'h4b9: dout <= -'sd28967; // 1209
        'h4ba: dout <= -'sd38818; // 1210
        'h4bb: dout <= -'sd42673; // 1211
        'h4bc: dout <= -'sd6454; // 1212
        'h4bd: dout <= -'sd53700; // 1213
        'h4be: dout <= -'sd46129; // 1214
        'h4bf: dout <= -'sd48466; // 1215
        'h4c0: dout <=  'sd13884; // 1216
        'h4c1: dout <=  'sd5322; // 1217
        'h4c2: dout <= -'sd34931; // 1218
        'h4c3: dout <= -'sd43208; // 1219
        'h4c4: dout <= -'sd48832; // 1220
        'h4c5: dout <=  'sd14947; // 1221
        'h4c6: dout <=  'sd36113; // 1222
        'h4c7: dout <=  'sd53909; // 1223
        'h4c8: dout <=  'sd56015; // 1224
        'h4c9: dout <= -'sd3916; // 1225
        'h4ca: dout <= -'sd44364; // 1226
        'h4cb: dout <= -'sd43102; // 1227
        'h4cc: dout <=  'sd8895; // 1228
        'h4cd: dout <= -'sd32272; // 1229
        'h4ce: dout <=  'sd6739; // 1230
        'h4cf: dout <= -'sd32071; // 1231
        'h4d0: dout <= -'sd36777; // 1232
        'h4d1: dout <=  'sd43771; // 1233
        'h4d2: dout <=  'sd14137; // 1234
        'h4d3: dout <=  'sd9152; // 1235
        'h4d4: dout <=  'sd1678; // 1236
        'h4d5: dout <=  'sd50531; // 1237
        'h4d6: dout <= -'sd32576; // 1238
        'h4d7: dout <= -'sd33883; // 1239
        'h4d8: dout <=  'sd2544; // 1240
        'h4d9: dout <= -'sd28982; // 1241
        'h4da: dout <=  'sd21799; // 1242
        'h4db: dout <= -'sd35668; // 1243
        'h4dc: dout <=  'sd32551; // 1244
        'h4dd: dout <= -'sd57111; // 1245
        'h4de: dout <= -'sd3623; // 1246
        'h4df: dout <=  'sd42649; // 1247
        'h4e0: dout <=  'sd4796; // 1248
        'h4e1: dout <= -'sd9623; // 1249
        'h4e2: dout <= -'sd260; // 1250
        'h4e3: dout <= -'sd43020; // 1251
        'h4e4: dout <=  'sd1888; // 1252
        'h4e5: dout <= -'sd48676; // 1253
        'h4e6: dout <=  'sd49678; // 1254
        'h4e7: dout <=  'sd8172; // 1255
        'h4e8: dout <= -'sd12469; // 1256
        'h4e9: dout <= -'sd9761; // 1257
        'h4ea: dout <= -'sd16695; // 1258
        'h4eb: dout <= -'sd48121; // 1259
        'h4ec: dout <=  'sd10060; // 1260
        'h4ed: dout <=  'sd7986; // 1261
        'h4ee: dout <= -'sd53447; // 1262
        'h4ef: dout <= -'sd27222; // 1263
        'h4f0: dout <=  'sd26645; // 1264
        'h4f1: dout <= -'sd53217; // 1265
        'h4f2: dout <=  'sd14157; // 1266
        'h4f3: dout <= -'sd1150; // 1267
        'h4f4: dout <=  'sd4387; // 1268
        'h4f5: dout <= -'sd24125; // 1269
        'h4f6: dout <= -'sd38647; // 1270
        'h4f7: dout <=  'sd14534; // 1271
        'h4f8: dout <=  'sd2822; // 1272
        'h4f9: dout <= -'sd18830; // 1273
        'h4fa: dout <=  'sd18445; // 1274
        'h4fb: dout <= -'sd1750; // 1275
        'h4fc: dout <=  'sd24398; // 1276
        'h4fd: dout <= -'sd39172; // 1277
        'h4fe: dout <=  'sd14131; // 1278
        'h4ff: dout <=  'sd49158; // 1279
        'h500: dout <=  'sd245; // 1280
        'h501: dout <= -'sd46560; // 1281
        'h502: dout <= -'sd41021; // 1282
        'h503: dout <=  'sd13573; // 1283
        'h504: dout <= -'sd15967; // 1284
        'h505: dout <= -'sd29372; // 1285
        'h506: dout <= -'sd42947; // 1286
        'h507: dout <= -'sd19152; // 1287
        'h508: dout <= -'sd54995; // 1288
        'h509: dout <= -'sd19960; // 1289
        'h50a: dout <=  'sd33234; // 1290
        'h50b: dout <= -'sd27099; // 1291
        'h50c: dout <= -'sd25473; // 1292
        'h50d: dout <= -'sd16934; // 1293
        'h50e: dout <= -'sd55098; // 1294
        'h50f: dout <=  'sd166; // 1295
        'h510: dout <=  'sd10569; // 1296
        'h511: dout <=  'sd21841; // 1297
        'h512: dout <=  'sd12931; // 1298
        'h513: dout <= -'sd22763; // 1299
        'h514: dout <= -'sd29479; // 1300
        'h515: dout <=  'sd5954; // 1301
        'h516: dout <=  'sd23950; // 1302
        'h517: dout <= -'sd10156; // 1303
        'h518: dout <=  'sd43868; // 1304
        'h519: dout <= -'sd29913; // 1305
        'h51a: dout <=  'sd33017; // 1306
        'h51b: dout <= -'sd18346; // 1307
        'h51c: dout <= -'sd54433; // 1308
        'h51d: dout <=  'sd30057; // 1309
        'h51e: dout <=  'sd14269; // 1310
        'h51f: dout <=  'sd44945; // 1311
        'h520: dout <= -'sd11928; // 1312
        'h521: dout <= -'sd51604; // 1313
        'h522: dout <= -'sd50209; // 1314
        'h523: dout <= -'sd14163; // 1315
        'h524: dout <=  'sd3172; // 1316
        'h525: dout <= -'sd24728; // 1317
        'h526: dout <=  'sd37888; // 1318
        'h527: dout <= -'sd1520; // 1319
        'h528: dout <= -'sd39082; // 1320
        'h529: dout <=  'sd16794; // 1321
        'h52a: dout <=  'sd8400; // 1322
        'h52b: dout <=  'sd52276; // 1323
        'h52c: dout <=  'sd5505; // 1324
        'h52d: dout <= -'sd27329; // 1325
        'h52e: dout <=  'sd49539; // 1326
        'h52f: dout <=  'sd25594; // 1327
        'h530: dout <=  'sd33351; // 1328
        'h531: dout <=  'sd18676; // 1329
        'h532: dout <= -'sd45410; // 1330
        'h533: dout <= -'sd15828; // 1331
        'h534: dout <= -'sd39577; // 1332
        'h535: dout <=  'sd36945; // 1333
        'h536: dout <= -'sd56965; // 1334
        'h537: dout <= -'sd22933; // 1335
        'h538: dout <= -'sd1786; // 1336
        'h539: dout <= -'sd3199; // 1337
        'h53a: dout <=  'sd14231; // 1338
        'h53b: dout <=  'sd27249; // 1339
        'h53c: dout <= -'sd639; // 1340
        'h53d: dout <= -'sd2107; // 1341
        'h53e: dout <=  'sd41728; // 1342
        'h53f: dout <= -'sd4125; // 1343
        'h540: dout <=  'sd26241; // 1344
        'h541: dout <=  'sd48726; // 1345
        'h542: dout <=  'sd51908; // 1346
        'h543: dout <=  'sd37068; // 1347
        'h544: dout <=  'sd44152; // 1348
        'h545: dout <= -'sd20593; // 1349
        'h546: dout <=  'sd45581; // 1350
        'h547: dout <= -'sd18491; // 1351
        'h548: dout <=  'sd9248; // 1352
        'h549: dout <= -'sd42108; // 1353
        'h54a: dout <=  'sd27773; // 1354
        'h54b: dout <= -'sd46414; // 1355
        'h54c: dout <=  'sd51227; // 1356
        'h54d: dout <= -'sd38186; // 1357
        'h54e: dout <=  'sd17524; // 1358
        'h54f: dout <= -'sd46377; // 1359
        'h550: dout <=  'sd52757; // 1360
        'h551: dout <= -'sd42572; // 1361
        'h552: dout <=  'sd27153; // 1362
        'h553: dout <= -'sd29569; // 1363
        'h554: dout <= -'sd44113; // 1364
        'h555: dout <= -'sd50676; // 1365
        'h556: dout <=  'sd33533; // 1366
        'h557: dout <= -'sd23262; // 1367
        'h558: dout <=  'sd31224; // 1368
        'h559: dout <=  'sd13983; // 1369
        'h55a: dout <= -'sd18437; // 1370
        'h55b: dout <=  'sd11927; // 1371
        'h55c: dout <=  'sd5815; // 1372
        'h55d: dout <= -'sd35935; // 1373
        'h55e: dout <=  'sd17046; // 1374
        'h55f: dout <= -'sd18393; // 1375
        'h560: dout <= -'sd16676; // 1376
        'h561: dout <= -'sd16170; // 1377
        'h562: dout <= -'sd22869; // 1378
        'h563: dout <= -'sd1171; // 1379
        'h564: dout <=  'sd43809; // 1380
        'h565: dout <=  'sd30918; // 1381
        'h566: dout <= -'sd8531; // 1382
        'h567: dout <=  'sd42166; // 1383
        'h568: dout <= -'sd14030; // 1384
        'h569: dout <= -'sd36684; // 1385
        'h56a: dout <= -'sd52978; // 1386
        'h56b: dout <=  'sd36344; // 1387
        'h56c: dout <=  'sd11688; // 1388
        'h56d: dout <=  'sd9200; // 1389
        'h56e: dout <= -'sd4382; // 1390
        'h56f: dout <= -'sd6172; // 1391
        'h570: dout <= -'sd48321; // 1392
        'h571: dout <=  'sd5436; // 1393
        'h572: dout <= -'sd43635; // 1394
        'h573: dout <=  'sd2710; // 1395
        'h574: dout <= -'sd40700; // 1396
        'h575: dout <= -'sd51513; // 1397
        'h576: dout <=  'sd19480; // 1398
        'h577: dout <=  'sd14608; // 1399
        'h578: dout <= -'sd31227; // 1400
        'h579: dout <= -'sd51870; // 1401
        'h57a: dout <= -'sd34531; // 1402
        'h57b: dout <= -'sd21839; // 1403
        'h57c: dout <= -'sd54216; // 1404
        'h57d: dout <= -'sd37730; // 1405
        'h57e: dout <= -'sd10355; // 1406
        'h57f: dout <= -'sd8952; // 1407
        'h580: dout <=  'sd14662; // 1408
        'h581: dout <= -'sd19064; // 1409
        'h582: dout <=  'sd8519; // 1410
        'h583: dout <=  'sd3231; // 1411
        'h584: dout <=  'sd20122; // 1412
        'h585: dout <= -'sd15673; // 1413
        'h586: dout <= -'sd8236; // 1414
        'h587: dout <= -'sd46138; // 1415
        'h588: dout <=  'sd23354; // 1416
        'h589: dout <= -'sd35375; // 1417
        'h58a: dout <=  'sd28742; // 1418
        'h58b: dout <=  'sd35051; // 1419
        'h58c: dout <= -'sd9961; // 1420
        'h58d: dout <= -'sd49397; // 1421
        'h58e: dout <=  'sd45256; // 1422
        'h58f: dout <= -'sd20033; // 1423
        'h590: dout <=  'sd10400; // 1424
        'h591: dout <= -'sd55698; // 1425
        'h592: dout <= -'sd13736; // 1426
        'h593: dout <=  'sd33424; // 1427
        'h594: dout <=  'sd51766; // 1428
        'h595: dout <=  'sd32982; // 1429
        'h596: dout <=  'sd17875; // 1430
        'h597: dout <=  'sd55354; // 1431
        'h598: dout <=  'sd32457; // 1432
        'h599: dout <=  'sd8074; // 1433
        'h59a: dout <=  'sd12645; // 1434
        'h59b: dout <= -'sd51017; // 1435
        'h59c: dout <= -'sd16708; // 1436
        'h59d: dout <=  'sd19018; // 1437
        'h59e: dout <=  'sd36248; // 1438
        'h59f: dout <=  'sd33565; // 1439
        'h5a0: dout <=  'sd14708; // 1440
        'h5a1: dout <= -'sd2839; // 1441
        'h5a2: dout <= -'sd14832; // 1442
        'h5a3: dout <=  'sd36489; // 1443
        'h5a4: dout <=  'sd46038; // 1444
        'h5a5: dout <= -'sd35013; // 1445
        'h5a6: dout <=  'sd6482; // 1446
        'h5a7: dout <= -'sd9978; // 1447
        'h5a8: dout <= -'sd7704; // 1448
        'h5a9: dout <=  'sd21723; // 1449
        'h5aa: dout <= -'sd36833; // 1450
        'h5ab: dout <= -'sd19334; // 1451
        'h5ac: dout <= -'sd6436; // 1452
        'h5ad: dout <= -'sd37953; // 1453
        'h5ae: dout <= -'sd9940; // 1454
        'h5af: dout <=  'sd29864; // 1455
        'h5b0: dout <= -'sd34671; // 1456
        'h5b1: dout <=  'sd25919; // 1457
        'h5b2: dout <=  'sd7345; // 1458
        'h5b3: dout <=  'sd1017; // 1459
        'h5b4: dout <=  'sd8412; // 1460
        'h5b5: dout <= -'sd53659; // 1461
        'h5b6: dout <=  'sd25847; // 1462
        'h5b7: dout <= -'sd23463; // 1463
        'h5b8: dout <= -'sd52386; // 1464
        'h5b9: dout <=  'sd46174; // 1465
        'h5ba: dout <= -'sd37506; // 1466
        'h5bb: dout <=  'sd20961; // 1467
        'h5bc: dout <= -'sd11404; // 1468
        'h5bd: dout <=  'sd17227; // 1469
        'h5be: dout <=  'sd16481; // 1470
        'h5bf: dout <= -'sd12327; // 1471
        'h5c0: dout <= -'sd51301; // 1472
        'h5c1: dout <= -'sd25388; // 1473
        'h5c2: dout <= -'sd20052; // 1474
        'h5c3: dout <= -'sd32306; // 1475
        'h5c4: dout <=  'sd5653; // 1476
        'h5c5: dout <=  'sd45804; // 1477
        'h5c6: dout <=  'sd21130; // 1478
        'h5c7: dout <=  'sd9511; // 1479
        'h5c8: dout <= -'sd46706; // 1480
        'h5c9: dout <=  'sd43372; // 1481
        'h5ca: dout <= -'sd11710; // 1482
        'h5cb: dout <=  'sd36218; // 1483
        'h5cc: dout <=  'sd22974; // 1484
        'h5cd: dout <= -'sd9309; // 1485
        'h5ce: dout <= -'sd35268; // 1486
        'h5cf: dout <= -'sd21480; // 1487
        'h5d0: dout <=  'sd20475; // 1488
        'h5d1: dout <=  'sd21057; // 1489
        'h5d2: dout <=  'sd30359; // 1490
        'h5d3: dout <=  'sd9826; // 1491
        'h5d4: dout <= -'sd46740; // 1492
        'h5d5: dout <= -'sd49304; // 1493
        'h5d6: dout <= -'sd1658; // 1494
        'h5d7: dout <= -'sd30103; // 1495
        'h5d8: dout <= -'sd24295; // 1496
        'h5d9: dout <=  'sd39455; // 1497
        'h5da: dout <= -'sd46302; // 1498
        'h5db: dout <=  'sd35880; // 1499
        'h5dc: dout <=  'sd23422; // 1500
        'h5dd: dout <=  'sd6800; // 1501
        'h5de: dout <=  'sd15411; // 1502
        'h5df: dout <= -'sd7669; // 1503
        'h5e0: dout <=  'sd36867; // 1504
        'h5e1: dout <= -'sd45688; // 1505
        'h5e2: dout <=  'sd50191; // 1506
        'h5e3: dout <=  'sd18322; // 1507
        'h5e4: dout <=  'sd7737; // 1508
        'h5e5: dout <= -'sd26590; // 1509
        'h5e6: dout <= -'sd39411; // 1510
        'h5e7: dout <=  'sd56319; // 1511
        'h5e8: dout <=  'sd19401; // 1512
        'h5e9: dout <=  'sd1632; // 1513
        'h5ea: dout <= -'sd1322; // 1514
        'h5eb: dout <= -'sd38246; // 1515
        'h5ec: dout <=  'sd26726; // 1516
        'h5ed: dout <= -'sd15795; // 1517
        'h5ee: dout <= -'sd18285; // 1518
        'h5ef: dout <=  'sd27320; // 1519
        'h5f0: dout <= -'sd54788; // 1520
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hq2_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [16:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'h000: dout <=  'sd33745; // 0
        'h001: dout <= -'sd30737; // 1
        'h002: dout <=  'sd27017; // 2
        'h003: dout <= -'sd49504; // 3
        'h004: dout <= -'sd31833; // 4
        'h005: dout <=  'sd2226; // 5
        'h006: dout <= -'sd3175; // 6
        'h007: dout <=  'sd8247; // 7
        'h008: dout <=  'sd7295; // 8
        'h009: dout <=  'sd34491; // 9
        'h00a: dout <= -'sd51817; // 10
        'h00b: dout <= -'sd40581; // 11
        'h00c: dout <=  'sd17497; // 12
        'h00d: dout <= -'sd49898; // 13
        'h00e: dout <= -'sd41442; // 14
        'h00f: dout <=  'sd58099; // 15
        'h010: dout <=  'sd47456; // 16
        'h011: dout <= -'sd57091; // 17
        'h012: dout <=  'sd6560; // 18
        'h013: dout <= -'sd41884; // 19
        'h014: dout <= -'sd34093; // 20
        'h015: dout <= -'sd27366; // 21
        'h016: dout <= -'sd10025; // 22
        'h017: dout <= -'sd38963; // 23
        'h018: dout <=  'sd60089; // 24
        'h019: dout <= -'sd58544; // 25
        'h01a: dout <=  'sd18255; // 26
        'h01b: dout <= -'sd12042; // 27
        'h01c: dout <=  'sd37284; // 28
        'h01d: dout <= -'sd9383; // 29
        'h01e: dout <=  'sd27067; // 30
        'h01f: dout <=  'sd45959; // 31
        'h020: dout <= -'sd54539; // 32
        'h021: dout <= -'sd45472; // 33
        'h022: dout <= -'sd17047; // 34
        'h023: dout <=  'sd4080; // 35
        'h024: dout <=  'sd36448; // 36
        'h025: dout <=  'sd915; // 37
        'h026: dout <= -'sd57422; // 38
        'h027: dout <=  'sd35490; // 39
        'h028: dout <=  'sd55081; // 40
        'h029: dout <=  'sd18183; // 41
        'h02a: dout <= -'sd38606; // 42
        'h02b: dout <=  'sd31854; // 43
        'h02c: dout <= -'sd1271; // 44
        'h02d: dout <=  'sd37378; // 45
        'h02e: dout <= -'sd49547; // 46
        'h02f: dout <= -'sd24033; // 47
        'h030: dout <= -'sd22983; // 48
        'h031: dout <= -'sd42433; // 49
        'h032: dout <= -'sd42511; // 50
        'h033: dout <= -'sd42973; // 51
        'h034: dout <=  'sd15815; // 52
        'h035: dout <=  'sd51181; // 53
        'h036: dout <=  'sd50728; // 54
        'h037: dout <= -'sd8332; // 55
        'h038: dout <=  'sd39007; // 56
        'h039: dout <=  'sd33218; // 57
        'h03a: dout <=  'sd52610; // 58
        'h03b: dout <=  'sd14755; // 59
        'h03c: dout <=  'sd24990; // 60
        'h03d: dout <=  'sd27881; // 61
        'h03e: dout <=  'sd4778; // 62
        'h03f: dout <= -'sd36397; // 63
        'h040: dout <=  'sd37608; // 64
        'h041: dout <=  'sd48286; // 65
        'h042: dout <= -'sd21463; // 66
        'h043: dout <= -'sd23866; // 67
        'h044: dout <= -'sd6594; // 68
        'h045: dout <=  'sd34855; // 69
        'h046: dout <= -'sd52328; // 70
        'h047: dout <= -'sd57538; // 71
        'h048: dout <=  'sd45913; // 72
        'h049: dout <= -'sd5261; // 73
        'h04a: dout <=  'sd30239; // 74
        'h04b: dout <=  'sd23481; // 75
        'h04c: dout <= -'sd9067; // 76
        'h04d: dout <= -'sd44284; // 77
        'h04e: dout <= -'sd50566; // 78
        'h04f: dout <=  'sd25839; // 79
        'h050: dout <=  'sd48138; // 80
        'h051: dout <= -'sd7439; // 81
        'h052: dout <= -'sd54434; // 82
        'h053: dout <=  'sd27124; // 83
        'h054: dout <= -'sd54479; // 84
        'h055: dout <=  'sd14741; // 85
        'h056: dout <= -'sd38047; // 86
        'h057: dout <= -'sd35721; // 87
        'h058: dout <= -'sd26159; // 88
        'h059: dout <=  'sd3414; // 89
        'h05a: dout <= -'sd56176; // 90
        'h05b: dout <= -'sd25400; // 91
        'h05c: dout <=  'sd183; // 92
        'h05d: dout <=  'sd49820; // 93
        'h05e: dout <=  'sd9726; // 94
        'h05f: dout <= -'sd5232; // 95
        'h060: dout <= -'sd37523; // 96
        'h061: dout <= -'sd2968; // 97
        'h062: dout <= -'sd29169; // 98
        'h063: dout <=  'sd18044; // 99
        'h064: dout <= -'sd11362; // 100
        'h065: dout <= -'sd57551; // 101
        'h066: dout <= -'sd44775; // 102
        'h067: dout <=  'sd57067; // 103
        'h068: dout <= -'sd6527; // 104
        'h069: dout <=  'sd11467; // 105
        'h06a: dout <=  'sd7536; // 106
        'h06b: dout <= -'sd47040; // 107
        'h06c: dout <=  'sd50881; // 108
        'h06d: dout <= -'sd28795; // 109
        'h06e: dout <= -'sd26051; // 110
        'h06f: dout <=  'sd38530; // 111
        'h070: dout <= -'sd27341; // 112
        'h071: dout <= -'sd49659; // 113
        'h072: dout <=  'sd37923; // 114
        'h073: dout <= -'sd30224; // 115
        'h074: dout <=  'sd28255; // 116
        'h075: dout <=  'sd7913; // 117
        'h076: dout <=  'sd14686; // 118
        'h077: dout <= -'sd1107; // 119
        'h078: dout <=  'sd4477; // 120
        'h079: dout <=  'sd33456; // 121
        'h07a: dout <=  'sd52578; // 122
        'h07b: dout <= -'sd9417; // 123
        'h07c: dout <=  'sd33939; // 124
        'h07d: dout <= -'sd52494; // 125
        'h07e: dout <= -'sd37721; // 126
        'h07f: dout <=  'sd16825; // 127
        'h080: dout <=  'sd34058; // 128
        'h081: dout <=  'sd34741; // 129
        'h082: dout <=  'sd9138; // 130
        'h083: dout <= -'sd53321; // 131
        'h084: dout <=  'sd33367; // 132
        'h085: dout <=  'sd22824; // 133
        'h086: dout <=  'sd6616; // 134
        'h087: dout <=  'sd26690; // 135
        'h088: dout <= -'sd18887; // 136
        'h089: dout <= -'sd38012; // 137
        'h08a: dout <= -'sd30098; // 138
        'h08b: dout <= -'sd30271; // 139
        'h08c: dout <= -'sd40681; // 140
        'h08d: dout <=  'sd27139; // 141
        'h08e: dout <= -'sd2945; // 142
        'h08f: dout <= -'sd28751; // 143
        'h090: dout <=  'sd46783; // 144
        'h091: dout <=  'sd31444; // 145
        'h092: dout <= -'sd14678; // 146
        'h093: dout <= -'sd24749; // 147
        'h094: dout <= -'sd47770; // 148
        'h095: dout <= -'sd31195; // 149
        'h096: dout <= -'sd55160; // 150
        'h097: dout <=  'sd14682; // 151
        'h098: dout <= -'sd1329; // 152
        'h099: dout <= -'sd35571; // 153
        'h09a: dout <=  'sd44007; // 154
        'h09b: dout <=  'sd58082; // 155
        'h09c: dout <=  'sd34325; // 156
        'h09d: dout <= -'sd14207; // 157
        'h09e: dout <= -'sd31884; // 158
        'h09f: dout <= -'sd42571; // 159
        'h0a0: dout <= -'sd3486; // 160
        'h0a1: dout <=  'sd31926; // 161
        'h0a2: dout <=  'sd20883; // 162
        'h0a3: dout <=  'sd54195; // 163
        'h0a4: dout <= -'sd6312; // 164
        'h0a5: dout <=  'sd43294; // 165
        'h0a6: dout <= -'sd56828; // 166
        'h0a7: dout <= -'sd17659; // 167
        'h0a8: dout <=  'sd8655; // 168
        'h0a9: dout <= -'sd14795; // 169
        'h0aa: dout <= -'sd9505; // 170
        'h0ab: dout <= -'sd37774; // 171
        'h0ac: dout <=  'sd1097; // 172
        'h0ad: dout <= -'sd28927; // 173
        'h0ae: dout <=  'sd57135; // 174
        'h0af: dout <= -'sd24031; // 175
        'h0b0: dout <= -'sd18627; // 176
        'h0b1: dout <=  'sd29778; // 177
        'h0b2: dout <= -'sd23486; // 178
        'h0b3: dout <= -'sd52970; // 179
        'h0b4: dout <=  'sd3410; // 180
        'h0b5: dout <=  'sd35236; // 181
        'h0b6: dout <=  'sd50554; // 182
        'h0b7: dout <= -'sd15501; // 183
        'h0b8: dout <=  'sd47121; // 184
        'h0b9: dout <= -'sd47322; // 185
        'h0ba: dout <= -'sd54341; // 186
        'h0bb: dout <= -'sd51863; // 187
        'h0bc: dout <= -'sd32142; // 188
        'h0bd: dout <=  'sd40206; // 189
        'h0be: dout <= -'sd34241; // 190
        'h0bf: dout <=  'sd43924; // 191
        'h0c0: dout <= -'sd18977; // 192
        'h0c1: dout <= -'sd2999; // 193
        'h0c2: dout <=  'sd37250; // 194
        'h0c3: dout <=  'sd9422; // 195
        'h0c4: dout <=  'sd32167; // 196
        'h0c5: dout <=  'sd25269; // 197
        'h0c6: dout <= -'sd32024; // 198
        'h0c7: dout <= -'sd55502; // 199
        'h0c8: dout <=  'sd26591; // 200
        'h0c9: dout <= -'sd13737; // 201
        'h0ca: dout <= -'sd15298; // 202
        'h0cb: dout <= -'sd24346; // 203
        'h0cc: dout <= -'sd24783; // 204
        'h0cd: dout <=  'sd29769; // 205
        'h0ce: dout <= -'sd22281; // 206
        'h0cf: dout <= -'sd37725; // 207
        'h0d0: dout <= -'sd21028; // 208
        'h0d1: dout <= -'sd25055; // 209
        'h0d2: dout <=  'sd12376; // 210
        'h0d3: dout <= -'sd21537; // 211
        'h0d4: dout <=  'sd47876; // 212
        'h0d5: dout <= -'sd8220; // 213
        'h0d6: dout <=  'sd58510; // 214
        'h0d7: dout <= -'sd30570; // 215
        'h0d8: dout <=  'sd55866; // 216
        'h0d9: dout <= -'sd45804; // 217
        'h0da: dout <= -'sd52536; // 218
        'h0db: dout <=  'sd38811; // 219
        'h0dc: dout <=  'sd56140; // 220
        'h0dd: dout <=  'sd27528; // 221
        'h0de: dout <=  'sd56125; // 222
        'h0df: dout <=  'sd21861; // 223
        'h0e0: dout <= -'sd32915; // 224
        'h0e1: dout <= -'sd15370; // 225
        'h0e2: dout <= -'sd2422; // 226
        'h0e3: dout <=  'sd46762; // 227
        'h0e4: dout <=  'sd10729; // 228
        'h0e5: dout <=  'sd48836; // 229
        'h0e6: dout <=  'sd11129; // 230
        'h0e7: dout <= -'sd10107; // 231
        'h0e8: dout <= -'sd1513; // 232
        'h0e9: dout <=  'sd59940; // 233
        'h0ea: dout <=  'sd32076; // 234
        'h0eb: dout <=  'sd5420; // 235
        'h0ec: dout <= -'sd14443; // 236
        'h0ed: dout <=  'sd31087; // 237
        'h0ee: dout <=  'sd52774; // 238
        'h0ef: dout <= -'sd14043; // 239
        'h0f0: dout <= -'sd59021; // 240
        'h0f1: dout <= -'sd4035; // 241
        'h0f2: dout <=  'sd38838; // 242
        'h0f3: dout <=  'sd13955; // 243
        'h0f4: dout <=  'sd15340; // 244
        'h0f5: dout <= -'sd33990; // 245
        'h0f6: dout <= -'sd19608; // 246
        'h0f7: dout <=  'sd57334; // 247
        'h0f8: dout <=  'sd12102; // 248
        'h0f9: dout <= -'sd58176; // 249
        'h0fa: dout <= -'sd55415; // 250
        'h0fb: dout <= -'sd32119; // 251
        'h0fc: dout <=  'sd46763; // 252
        'h0fd: dout <=  'sd26094; // 253
        'h0fe: dout <= -'sd17437; // 254
        'h0ff: dout <=  'sd22352; // 255
        'h100: dout <=  'sd38914; // 256
        'h101: dout <= -'sd56019; // 257
        'h102: dout <=  'sd2656; // 258
        'h103: dout <=  'sd20252; // 259
        'h104: dout <= -'sd6070; // 260
        'h105: dout <=  'sd56123; // 261
        'h106: dout <= -'sd13661; // 262
        'h107: dout <=  'sd48573; // 263
        'h108: dout <= -'sd6139; // 264
        'h109: dout <= -'sd35950; // 265
        'h10a: dout <=  'sd9479; // 266
        'h10b: dout <=  'sd20771; // 267
        'h10c: dout <=  'sd21754; // 268
        'h10d: dout <= -'sd43506; // 269
        'h10e: dout <= -'sd52406; // 270
        'h10f: dout <= -'sd40875; // 271
        'h110: dout <=  'sd10938; // 272
        'h111: dout <= -'sd43392; // 273
        'h112: dout <= -'sd14165; // 274
        'h113: dout <= -'sd33763; // 275
        'h114: dout <= -'sd35168; // 276
        'h115: dout <= -'sd26144; // 277
        'h116: dout <=  'sd37911; // 278
        'h117: dout <= -'sd15992; // 279
        'h118: dout <=  'sd58435; // 280
        'h119: dout <= -'sd9109; // 281
        'h11a: dout <= -'sd50760; // 282
        'h11b: dout <=  'sd17746; // 283
        'h11c: dout <= -'sd36708; // 284
        'h11d: dout <= -'sd18398; // 285
        'h11e: dout <= -'sd7530; // 286
        'h11f: dout <=  'sd18257; // 287
        'h120: dout <=  'sd56050; // 288
        'h121: dout <= -'sd823; // 289
        'h122: dout <= -'sd12583; // 290
        'h123: dout <=  'sd58156; // 291
        'h124: dout <=  'sd25839; // 292
        'h125: dout <= -'sd50253; // 293
        'h126: dout <= -'sd59245; // 294
        'h127: dout <= -'sd7224; // 295
        'h128: dout <= -'sd6746; // 296
        'h129: dout <=  'sd31584; // 297
        'h12a: dout <= -'sd52702; // 298
        'h12b: dout <= -'sd46439; // 299
        'h12c: dout <=  'sd56904; // 300
        'h12d: dout <= -'sd26290; // 301
        'h12e: dout <=  'sd21696; // 302
        'h12f: dout <=  'sd52273; // 303
        'h130: dout <= -'sd13353; // 304
        'h131: dout <= -'sd46044; // 305
        'h132: dout <=  'sd5182; // 306
        'h133: dout <=  'sd22881; // 307
        'h134: dout <=  'sd11919; // 308
        'h135: dout <=  'sd13360; // 309
        'h136: dout <=  'sd51116; // 310
        'h137: dout <=  'sd48129; // 311
        'h138: dout <= -'sd39612; // 312
        'h139: dout <=  'sd48258; // 313
        'h13a: dout <=  'sd51721; // 314
        'h13b: dout <= -'sd30124; // 315
        'h13c: dout <= -'sd4676; // 316
        'h13d: dout <=  'sd8021; // 317
        'h13e: dout <=  'sd47429; // 318
        'h13f: dout <=  'sd52246; // 319
        'h140: dout <= -'sd16148; // 320
        'h141: dout <=  'sd43892; // 321
        'h142: dout <= -'sd33892; // 322
        'h143: dout <=  'sd1481; // 323
        'h144: dout <=  'sd20652; // 324
        'h145: dout <=  'sd15305; // 325
        'h146: dout <= -'sd38071; // 326
        'h147: dout <= -'sd35453; // 327
        'h148: dout <=  'sd39536; // 328
        'h149: dout <= -'sd59017; // 329
        'h14a: dout <=  'sd33038; // 330
        'h14b: dout <=  'sd46195; // 331
        'h14c: dout <= -'sd25085; // 332
        'h14d: dout <=  'sd55491; // 333
        'h14e: dout <= -'sd5341; // 334
        'h14f: dout <=  'sd46856; // 335
        'h150: dout <= -'sd9119; // 336
        'h151: dout <= -'sd56523; // 337
        'h152: dout <=  'sd20271; // 338
        'h153: dout <=  'sd48250; // 339
        'h154: dout <=  'sd53407; // 340
        'h155: dout <= -'sd17075; // 341
        'h156: dout <=  'sd34107; // 342
        'h157: dout <=  'sd1400; // 343
        'h158: dout <=  'sd22413; // 344
        'h159: dout <= -'sd18043; // 345
        'h15a: dout <=  'sd5516; // 346
        'h15b: dout <=  'sd48697; // 347
        'h15c: dout <=  'sd14264; // 348
        'h15d: dout <=  'sd45099; // 349
        'h15e: dout <= -'sd46543; // 350
        'h15f: dout <=  'sd26199; // 351
        'h160: dout <=  'sd8613; // 352
        'h161: dout <= -'sd7002; // 353
        'h162: dout <=  'sd54448; // 354
        'h163: dout <=  'sd48992; // 355
        'h164: dout <=  'sd1900; // 356
        'h165: dout <=  'sd16951; // 357
        'h166: dout <=  'sd54180; // 358
        'h167: dout <= -'sd46303; // 359
        'h168: dout <= -'sd57455; // 360
        'h169: dout <=  'sd49038; // 361
        'h16a: dout <= -'sd18661; // 362
        'h16b: dout <= -'sd48804; // 363
        'h16c: dout <=  'sd2738; // 364
        'h16d: dout <=  'sd145; // 365
        'h16e: dout <=  'sd53566; // 366
        'h16f: dout <= -'sd17399; // 367
        'h170: dout <=  'sd14048; // 368
        'h171: dout <=  'sd45313; // 369
        'h172: dout <=  'sd27152; // 370
        'h173: dout <=  'sd46284; // 371
        'h174: dout <=  'sd5597; // 372
        'h175: dout <=  'sd8183; // 373
        'h176: dout <= -'sd41762; // 374
        'h177: dout <=  'sd5167; // 375
        'h178: dout <=  'sd48123; // 376
        'h179: dout <= -'sd48767; // 377
        'h17a: dout <= -'sd42775; // 378
        'h17b: dout <=  'sd57891; // 379
        'h17c: dout <= -'sd51206; // 380
        'h17d: dout <=  'sd42295; // 381
        'h17e: dout <=  'sd40744; // 382
        'h17f: dout <=  'sd50327; // 383
        'h180: dout <= -'sd55596; // 384
        'h181: dout <=  'sd30018; // 385
        'h182: dout <= -'sd47358; // 386
        'h183: dout <= -'sd40816; // 387
        'h184: dout <=  'sd47419; // 388
        'h185: dout <=  'sd8967; // 389
        'h186: dout <=  'sd44565; // 390
        'h187: dout <=  'sd27285; // 391
        'h188: dout <=  'sd51582; // 392
        'h189: dout <= -'sd8285; // 393
        'h18a: dout <=  'sd5513; // 394
        'h18b: dout <= -'sd46027; // 395
        'h18c: dout <=  'sd387; // 396
        'h18d: dout <= -'sd19624; // 397
        'h18e: dout <=  'sd21931; // 398
        'h18f: dout <= -'sd18827; // 399
        'h190: dout <= -'sd46573; // 400
        'h191: dout <=  'sd41168; // 401
        'h192: dout <=  'sd49075; // 402
        'h193: dout <= -'sd46304; // 403
        'h194: dout <=  'sd47863; // 404
        'h195: dout <=  'sd29816; // 405
        'h196: dout <=  'sd51060; // 406
        'h197: dout <= -'sd47208; // 407
        'h198: dout <=  'sd40989; // 408
        'h199: dout <=  'sd45114; // 409
        'h19a: dout <= -'sd14690; // 410
        'h19b: dout <=  'sd24636; // 411
        'h19c: dout <=  'sd53965; // 412
        'h19d: dout <=  'sd2323; // 413
        'h19e: dout <= -'sd17630; // 414
        'h19f: dout <=  'sd50283; // 415
        'h1a0: dout <=  'sd29038; // 416
        'h1a1: dout <=  'sd37262; // 417
        'h1a2: dout <= -'sd11724; // 418
        'h1a3: dout <= -'sd35973; // 419
        'h1a4: dout <= -'sd46900; // 420
        'h1a5: dout <= -'sd22095; // 421
        'h1a6: dout <=  'sd5655; // 422
        'h1a7: dout <= -'sd31613; // 423
        'h1a8: dout <=  'sd13894; // 424
        'h1a9: dout <=  'sd21906; // 425
        'h1aa: dout <= -'sd10522; // 426
        'h1ab: dout <= -'sd45455; // 427
        'h1ac: dout <=  'sd9616; // 428
        'h1ad: dout <=  'sd39937; // 429
        'h1ae: dout <=  'sd41442; // 430
        'h1af: dout <=  'sd7104; // 431
        'h1b0: dout <= -'sd52036; // 432
        'h1b1: dout <= -'sd27109; // 433
        'h1b2: dout <=  'sd42562; // 434
        'h1b3: dout <= -'sd55957; // 435
        'h1b4: dout <=  'sd20066; // 436
        'h1b5: dout <= -'sd2324; // 437
        'h1b6: dout <=  'sd36627; // 438
        'h1b7: dout <=  'sd59064; // 439
        'h1b8: dout <= -'sd39361; // 440
        'h1b9: dout <= -'sd45745; // 441
        'h1ba: dout <=  'sd37900; // 442
        'h1bb: dout <= -'sd2512; // 443
        'h1bc: dout <=  'sd15271; // 444
        'h1bd: dout <= -'sd22989; // 445
        'h1be: dout <=  'sd18991; // 446
        'h1bf: dout <= -'sd19952; // 447
        'h1c0: dout <=  'sd14682; // 448
        'h1c1: dout <= -'sd47930; // 449
        'h1c2: dout <= -'sd48166; // 450
        'h1c3: dout <= -'sd32518; // 451
        'h1c4: dout <= -'sd49558; // 452
        'h1c5: dout <= -'sd48357; // 453
        'h1c6: dout <=  'sd53123; // 454
        'h1c7: dout <= -'sd16324; // 455
        'h1c8: dout <=  'sd28675; // 456
        'h1c9: dout <= -'sd22048; // 457
        'h1ca: dout <=  'sd9415; // 458
        'h1cb: dout <= -'sd11424; // 459
        'h1cc: dout <=  'sd18882; // 460
        'h1cd: dout <= -'sd28021; // 461
        'h1ce: dout <=  'sd30118; // 462
        'h1cf: dout <=  'sd39193; // 463
        'h1d0: dout <=  'sd17828; // 464
        'h1d1: dout <=  'sd26414; // 465
        'h1d2: dout <= -'sd35439; // 466
        'h1d3: dout <= -'sd60325; // 467
        'h1d4: dout <= -'sd39143; // 468
        'h1d5: dout <=  'sd47941; // 469
        'h1d6: dout <= -'sd17917; // 470
        'h1d7: dout <=  'sd1291; // 471
        'h1d8: dout <= -'sd33681; // 472
        'h1d9: dout <=  'sd30043; // 473
        'h1da: dout <= -'sd18580; // 474
        'h1db: dout <=  'sd38430; // 475
        'h1dc: dout <= -'sd49750; // 476
        'h1dd: dout <=  'sd44627; // 477
        'h1de: dout <= -'sd23660; // 478
        'h1df: dout <= -'sd48207; // 479
        'h1e0: dout <= -'sd16579; // 480
        'h1e1: dout <= -'sd25509; // 481
        'h1e2: dout <=  'sd58808; // 482
        'h1e3: dout <=  'sd22461; // 483
        'h1e4: dout <= -'sd2233; // 484
        'h1e5: dout <= -'sd292; // 485
        'h1e6: dout <= -'sd20016; // 486
        'h1e7: dout <= -'sd58725; // 487
        'h1e8: dout <=  'sd43607; // 488
        'h1e9: dout <= -'sd10009; // 489
        'h1ea: dout <= -'sd4688; // 490
        'h1eb: dout <= -'sd30264; // 491
        'h1ec: dout <=  'sd37164; // 492
        'h1ed: dout <= -'sd44494; // 493
        'h1ee: dout <= -'sd22048; // 494
        'h1ef: dout <= -'sd34567; // 495
        'h1f0: dout <= -'sd16949; // 496
        'h1f1: dout <=  'sd33801; // 497
        'h1f2: dout <= -'sd22988; // 498
        'h1f3: dout <= -'sd36534; // 499
        'h1f4: dout <=  'sd39705; // 500
        'h1f5: dout <=  'sd45635; // 501
        'h1f6: dout <=  'sd31266; // 502
        'h1f7: dout <=  'sd7969; // 503
        'h1f8: dout <= -'sd34526; // 504
        'h1f9: dout <=  'sd16037; // 505
        'h1fa: dout <=  'sd16295; // 506
        'h1fb: dout <= -'sd43169; // 507
        'h1fc: dout <= -'sd44014; // 508
        'h1fd: dout <=  'sd8241; // 509
        'h1fe: dout <= -'sd52079; // 510
        'h1ff: dout <=  'sd1084; // 511
        'h200: dout <=  'sd30390; // 512
        'h201: dout <=  'sd29517; // 513
        'h202: dout <= -'sd7594; // 514
        'h203: dout <= -'sd51607; // 515
        'h204: dout <= -'sd12479; // 516
        'h205: dout <=  'sd40991; // 517
        'h206: dout <= -'sd60300; // 518
        'h207: dout <= -'sd36235; // 519
        'h208: dout <= -'sd43732; // 520
        'h209: dout <= -'sd20140; // 521
        'h20a: dout <= -'sd60247; // 522
        'h20b: dout <=  'sd6131; // 523
        'h20c: dout <= -'sd59308; // 524
        'h20d: dout <=  'sd22582; // 525
        'h20e: dout <=  'sd449; // 526
        'h20f: dout <=  'sd28213; // 527
        'h210: dout <=  'sd24007; // 528
        'h211: dout <= -'sd40470; // 529
        'h212: dout <=  'sd48487; // 530
        'h213: dout <=  'sd14168; // 531
        'h214: dout <=  'sd31223; // 532
        'h215: dout <= -'sd42207; // 533
        'h216: dout <= -'sd58542; // 534
        'h217: dout <= -'sd19459; // 535
        'h218: dout <=  'sd33429; // 536
        'h219: dout <= -'sd30621; // 537
        'h21a: dout <= -'sd26536; // 538
        'h21b: dout <=  'sd53353; // 539
        'h21c: dout <=  'sd59214; // 540
        'h21d: dout <=  'sd36312; // 541
        'h21e: dout <= -'sd30225; // 542
        'h21f: dout <= -'sd32104; // 543
        'h220: dout <=  'sd60399; // 544
        'h221: dout <=  'sd47753; // 545
        'h222: dout <= -'sd35391; // 546
        'h223: dout <= -'sd18648; // 547
        'h224: dout <= -'sd16904; // 548
        'h225: dout <=  'sd36992; // 549
        'h226: dout <=  'sd23485; // 550
        'h227: dout <= -'sd43855; // 551
        'h228: dout <= -'sd55577; // 552
        'h229: dout <=  'sd13341; // 553
        'h22a: dout <=  'sd6445; // 554
        'h22b: dout <=  'sd56257; // 555
        'h22c: dout <=  'sd46229; // 556
        'h22d: dout <=  'sd23145; // 557
        'h22e: dout <= -'sd38326; // 558
        'h22f: dout <= -'sd12113; // 559
        'h230: dout <= -'sd35793; // 560
        'h231: dout <= -'sd681; // 561
        'h232: dout <=  'sd20985; // 562
        'h233: dout <=  'sd35764; // 563
        'h234: dout <=  'sd7563; // 564
        'h235: dout <= -'sd14055; // 565
        'h236: dout <=  'sd5983; // 566
        'h237: dout <= -'sd49366; // 567
        'h238: dout <=  'sd646; // 568
        'h239: dout <= -'sd51885; // 569
        'h23a: dout <= -'sd56689; // 570
        'h23b: dout <= -'sd17012; // 571
        'h23c: dout <= -'sd483; // 572
        'h23d: dout <= -'sd19435; // 573
        'h23e: dout <=  'sd59686; // 574
        'h23f: dout <=  'sd48435; // 575
        'h240: dout <=  'sd18816; // 576
        'h241: dout <= -'sd27153; // 577
        'h242: dout <=  'sd52890; // 578
        'h243: dout <=  'sd10556; // 579
        'h244: dout <= -'sd50557; // 580
        'h245: dout <= -'sd51018; // 581
        'h246: dout <= -'sd13972; // 582
        'h247: dout <=  'sd46582; // 583
        'h248: dout <= -'sd48009; // 584
        'h249: dout <=  'sd58809; // 585
        'h24a: dout <=  'sd12333; // 586
        'h24b: dout <=  'sd57126; // 587
        'h24c: dout <=  'sd36282; // 588
        'h24d: dout <=  'sd34102; // 589
        'h24e: dout <=  'sd9624; // 590
        'h24f: dout <= -'sd40611; // 591
        'h250: dout <= -'sd30694; // 592
        'h251: dout <= -'sd41551; // 593
        'h252: dout <=  'sd39849; // 594
        'h253: dout <=  'sd6534; // 595
        'h254: dout <=  'sd17964; // 596
        'h255: dout <= -'sd3835; // 597
        'h256: dout <=  'sd16958; // 598
        'h257: dout <= -'sd14568; // 599
        'h258: dout <=  'sd2598; // 600
        'h259: dout <= -'sd38456; // 601
        'h25a: dout <= -'sd55955; // 602
        'h25b: dout <= -'sd34658; // 603
        'h25c: dout <= -'sd52043; // 604
        'h25d: dout <= -'sd35181; // 605
        'h25e: dout <= -'sd55825; // 606
        'h25f: dout <= -'sd2034; // 607
        'h260: dout <=  'sd56864; // 608
        'h261: dout <=  'sd8918; // 609
        'h262: dout <=  'sd49906; // 610
        'h263: dout <= -'sd35477; // 611
        'h264: dout <=  'sd12202; // 612
        'h265: dout <=  'sd29029; // 613
        'h266: dout <=  'sd8172; // 614
        'h267: dout <=  'sd15201; // 615
        'h268: dout <=  'sd41803; // 616
        'h269: dout <=  'sd23463; // 617
        'h26a: dout <=  'sd53686; // 618
        'h26b: dout <= -'sd56645; // 619
        'h26c: dout <=  'sd37212; // 620
        'h26d: dout <=  'sd26569; // 621
        'h26e: dout <= -'sd13150; // 622
        'h26f: dout <= -'sd59136; // 623
        'h270: dout <= -'sd23089; // 624
        'h271: dout <= -'sd36681; // 625
        'h272: dout <= -'sd30549; // 626
        'h273: dout <= -'sd35612; // 627
        'h274: dout <=  'sd48608; // 628
        'h275: dout <= -'sd3736; // 629
        'h276: dout <=  'sd29409; // 630
        'h277: dout <=  'sd58612; // 631
        'h278: dout <=  'sd41499; // 632
        'h279: dout <= -'sd46706; // 633
        'h27a: dout <= -'sd28974; // 634
        'h27b: dout <= -'sd3015; // 635
        'h27c: dout <=  'sd27173; // 636
        'h27d: dout <=  'sd48533; // 637
        'h27e: dout <=  'sd44473; // 638
        'h27f: dout <=  'sd14906; // 639
        'h280: dout <=  'sd53029; // 640
        'h281: dout <=  'sd49662; // 641
        'h282: dout <= -'sd34464; // 642
        'h283: dout <=  'sd6753; // 643
        'h284: dout <=  'sd5956; // 644
        'h285: dout <=  'sd42745; // 645
        'h286: dout <= -'sd50453; // 646
        'h287: dout <=  'sd4625; // 647
        'h288: dout <=  'sd33070; // 648
        'h289: dout <=  'sd31489; // 649
        'h28a: dout <= -'sd15756; // 650
        'h28b: dout <= -'sd31133; // 651
        'h28c: dout <=  'sd53494; // 652
        'h28d: dout <= -'sd37543; // 653
        'h28e: dout <= -'sd54020; // 654
        'h28f: dout <= -'sd49314; // 655
        'h290: dout <=  'sd13178; // 656
        'h291: dout <= -'sd54981; // 657
        'h292: dout <=  'sd11346; // 658
        'h293: dout <= -'sd16371; // 659
        'h294: dout <= -'sd8830; // 660
        'h295: dout <=  'sd22979; // 661
        'h296: dout <=  'sd35032; // 662
        'h297: dout <= -'sd16240; // 663
        'h298: dout <= -'sd21475; // 664
        'h299: dout <= -'sd5928; // 665
        'h29a: dout <=  'sd28087; // 666
        'h29b: dout <= -'sd16611; // 667
        'h29c: dout <= -'sd38685; // 668
        'h29d: dout <= -'sd17452; // 669
        'h29e: dout <=  'sd8525; // 670
        'h29f: dout <=  'sd10852; // 671
        'h2a0: dout <= -'sd24803; // 672
        'h2a1: dout <=  'sd22020; // 673
        'h2a2: dout <=  'sd8420; // 674
        'h2a3: dout <= -'sd32130; // 675
        'h2a4: dout <= -'sd3496; // 676
        'h2a5: dout <= -'sd20145; // 677
        'h2a6: dout <=  'sd20910; // 678
        'h2a7: dout <= -'sd39577; // 679
        'h2a8: dout <= -'sd54755; // 680
        'h2a9: dout <= -'sd10841; // 681
        'h2aa: dout <= -'sd30475; // 682
        'h2ab: dout <= -'sd8813; // 683
        'h2ac: dout <= -'sd54787; // 684
        'h2ad: dout <=  'sd58452; // 685
        'h2ae: dout <= -'sd53261; // 686
        'h2af: dout <=  'sd28382; // 687
        'h2b0: dout <=  'sd3884; // 688
        'h2b1: dout <=  'sd21217; // 689
        'h2b2: dout <= -'sd59011; // 690
        'h2b3: dout <= -'sd48799; // 691
        'h2b4: dout <=  'sd40066; // 692
        'h2b5: dout <=  'sd27643; // 693
        'h2b6: dout <=  'sd33223; // 694
        'h2b7: dout <=  'sd8610; // 695
        'h2b8: dout <=  'sd12865; // 696
        'h2b9: dout <= -'sd10773; // 697
        'h2ba: dout <= -'sd43611; // 698
        'h2bb: dout <= -'sd18155; // 699
        'h2bc: dout <= -'sd33670; // 700
        'h2bd: dout <=  'sd55646; // 701
        'h2be: dout <=  'sd45402; // 702
        'h2bf: dout <=  'sd771; // 703
        'h2c0: dout <= -'sd40907; // 704
        'h2c1: dout <=  'sd60353; // 705
        'h2c2: dout <= -'sd10843; // 706
        'h2c3: dout <= -'sd42657; // 707
        'h2c4: dout <= -'sd47035; // 708
        'h2c5: dout <= -'sd58496; // 709
        'h2c6: dout <=  'sd11672; // 710
        'h2c7: dout <=  'sd48164; // 711
        'h2c8: dout <= -'sd16725; // 712
        'h2c9: dout <= -'sd8699; // 713
        'h2ca: dout <=  'sd30343; // 714
        'h2cb: dout <=  'sd41630; // 715
        'h2cc: dout <= -'sd31767; // 716
        'h2cd: dout <=  'sd3630; // 717
        'h2ce: dout <=  'sd22454; // 718
        'h2cf: dout <= -'sd5357; // 719
        'h2d0: dout <=  'sd16604; // 720
        'h2d1: dout <=  'sd46324; // 721
        'h2d2: dout <=  'sd256; // 722
        'h2d3: dout <= -'sd13467; // 723
        'h2d4: dout <= -'sd24028; // 724
        'h2d5: dout <= -'sd13580; // 725
        'h2d6: dout <=  'sd16816; // 726
        'h2d7: dout <= -'sd9335; // 727
        'h2d8: dout <= -'sd45855; // 728
        'h2d9: dout <= -'sd45521; // 729
        'h2da: dout <=  'sd11893; // 730
        'h2db: dout <= -'sd30011; // 731
        'h2dc: dout <=  'sd9882; // 732
        'h2dd: dout <=  'sd37643; // 733
        'h2de: dout <=  'sd31119; // 734
        'h2df: dout <=  'sd37435; // 735
        'h2e0: dout <= -'sd53993; // 736
        'h2e1: dout <= -'sd9218; // 737
        'h2e2: dout <=  'sd35912; // 738
        'h2e3: dout <= -'sd20778; // 739
        'h2e4: dout <=  'sd50819; // 740
        'h2e5: dout <=  'sd14194; // 741
        'h2e6: dout <=  'sd52308; // 742
        'h2e7: dout <=  'sd29035; // 743
        'h2e8: dout <=  'sd31114; // 744
        'h2e9: dout <= -'sd41717; // 745
        'h2ea: dout <=  'sd55865; // 746
        'h2eb: dout <=  'sd7511; // 747
        'h2ec: dout <= -'sd10529; // 748
        'h2ed: dout <=  'sd49130; // 749
        'h2ee: dout <= -'sd38697; // 750
        'h2ef: dout <= -'sd33858; // 751
        'h2f0: dout <= -'sd47302; // 752
        'h2f1: dout <=  'sd53488; // 753
        'h2f2: dout <= -'sd48794; // 754
        'h2f3: dout <=  'sd598; // 755
        'h2f4: dout <=  'sd6403; // 756
        'h2f5: dout <= -'sd58971; // 757
        'h2f6: dout <=  'sd39521; // 758
        'h2f7: dout <= -'sd10187; // 759
        'h2f8: dout <=  'sd2409; // 760
        'h2f9: dout <= -'sd24900; // 761
        'h2fa: dout <= -'sd44797; // 762
        'h2fb: dout <= -'sd11730; // 763
        'h2fc: dout <= -'sd52330; // 764
        'h2fd: dout <= -'sd5155; // 765
        'h2fe: dout <=  'sd30009; // 766
        'h2ff: dout <= -'sd845; // 767
        'h300: dout <=  'sd54332; // 768
        'h301: dout <=  'sd30931; // 769
        'h302: dout <=  'sd37148; // 770
        'h303: dout <=  'sd41674; // 771
        'h304: dout <= -'sd11181; // 772
        'h305: dout <=  'sd41821; // 773
        'h306: dout <= -'sd5226; // 774
        'h307: dout <= -'sd30098; // 775
        'h308: dout <= -'sd12502; // 776
        'h309: dout <= -'sd54848; // 777
        'h30a: dout <=  'sd60039; // 778
        'h30b: dout <= -'sd42304; // 779
        'h30c: dout <=  'sd58203; // 780
        'h30d: dout <= -'sd22355; // 781
        'h30e: dout <=  'sd14766; // 782
        'h30f: dout <=  'sd53174; // 783
        'h310: dout <=  'sd38209; // 784
        'h311: dout <= -'sd42732; // 785
        'h312: dout <= -'sd31035; // 786
        'h313: dout <=  'sd10219; // 787
        'h314: dout <=  'sd52337; // 788
        'h315: dout <=  'sd11287; // 789
        'h316: dout <= -'sd15252; // 790
        'h317: dout <= -'sd49018; // 791
        'h318: dout <=  'sd5235; // 792
        'h319: dout <=  'sd17822; // 793
        'h31a: dout <=  'sd31049; // 794
        'h31b: dout <= -'sd30664; // 795
        'h31c: dout <= -'sd46272; // 796
        'h31d: dout <=  'sd54880; // 797
        'h31e: dout <= -'sd271; // 798
        'h31f: dout <= -'sd3354; // 799
        'h320: dout <= -'sd27192; // 800
        'h321: dout <= -'sd27350; // 801
        'h322: dout <=  'sd25603; // 802
        'h323: dout <=  'sd17025; // 803
        'h324: dout <=  'sd44813; // 804
        'h325: dout <=  'sd13756; // 805
        'h326: dout <= -'sd46427; // 806
        'h327: dout <=  'sd11162; // 807
        'h328: dout <=  'sd15072; // 808
        'h329: dout <=  'sd59688; // 809
        'h32a: dout <= -'sd763; // 810
        'h32b: dout <= -'sd30349; // 811
        'h32c: dout <=  'sd55916; // 812
        'h32d: dout <=  'sd36342; // 813
        'h32e: dout <= -'sd9174; // 814
        'h32f: dout <=  'sd57923; // 815
        'h330: dout <= -'sd10689; // 816
        'h331: dout <=  'sd19140; // 817
        'h332: dout <= -'sd9932; // 818
        'h333: dout <= -'sd16601; // 819
        'h334: dout <= -'sd24814; // 820
        'h335: dout <= -'sd48314; // 821
        'h336: dout <= -'sd54869; // 822
        'h337: dout <= -'sd56795; // 823
        'h338: dout <= -'sd35822; // 824
        'h339: dout <= -'sd2324; // 825
        'h33a: dout <= -'sd39558; // 826
        'h33b: dout <=  'sd12426; // 827
        'h33c: dout <=  'sd38410; // 828
        'h33d: dout <= -'sd46296; // 829
        'h33e: dout <=  'sd35717; // 830
        'h33f: dout <= -'sd53468; // 831
        'h340: dout <= -'sd41444; // 832
        'h341: dout <= -'sd53464; // 833
        'h342: dout <=  'sd58938; // 834
        'h343: dout <= -'sd24125; // 835
        'h344: dout <=  'sd29723; // 836
        'h345: dout <=  'sd50666; // 837
        'h346: dout <= -'sd15860; // 838
        'h347: dout <= -'sd19171; // 839
        'h348: dout <=  'sd7286; // 840
        'h349: dout <=  'sd55484; // 841
        'h34a: dout <= -'sd47278; // 842
        'h34b: dout <= -'sd59725; // 843
        'h34c: dout <= -'sd41409; // 844
        'h34d: dout <=  'sd48225; // 845
        'h34e: dout <= -'sd35691; // 846
        'h34f: dout <= -'sd14821; // 847
        'h350: dout <=  'sd28940; // 848
        'h351: dout <= -'sd34739; // 849
        'h352: dout <=  'sd58521; // 850
        'h353: dout <=  'sd46368; // 851
        'h354: dout <= -'sd41003; // 852
        'h355: dout <=  'sd57777; // 853
        'h356: dout <= -'sd4365; // 854
        'h357: dout <= -'sd31743; // 855
        'h358: dout <= -'sd11007; // 856
        'h359: dout <=  'sd11984; // 857
        'h35a: dout <= -'sd37306; // 858
        'h35b: dout <= -'sd14380; // 859
        'h35c: dout <=  'sd23855; // 860
        'h35d: dout <=  'sd21864; // 861
        'h35e: dout <=  'sd20876; // 862
        'h35f: dout <= -'sd17364; // 863
        'h360: dout <=  'sd8514; // 864
        'h361: dout <= -'sd26683; // 865
        'h362: dout <= -'sd32373; // 866
        'h363: dout <=  'sd38878; // 867
        'h364: dout <= -'sd2585; // 868
        'h365: dout <=  'sd42507; // 869
        'h366: dout <=  'sd54433; // 870
        'h367: dout <=  'sd32434; // 871
        'h368: dout <=  'sd28365; // 872
        'h369: dout <= -'sd53164; // 873
        'h36a: dout <= -'sd4477; // 874
        'h36b: dout <= -'sd24236; // 875
        'h36c: dout <=  'sd54483; // 876
        'h36d: dout <=  'sd12980; // 877
        'h36e: dout <=  'sd29188; // 878
        'h36f: dout <= -'sd49161; // 879
        'h370: dout <=  'sd14895; // 880
        'h371: dout <=  'sd23970; // 881
        'h372: dout <=  'sd11354; // 882
        'h373: dout <=  'sd24354; // 883
        'h374: dout <= -'sd2403; // 884
        'h375: dout <=  'sd7604; // 885
        'h376: dout <= -'sd1458; // 886
        'h377: dout <= -'sd7395; // 887
        'h378: dout <= -'sd34252; // 888
        'h379: dout <= -'sd15420; // 889
        'h37a: dout <=  'sd43642; // 890
        'h37b: dout <=  'sd42578; // 891
        'h37c: dout <=  'sd36135; // 892
        'h37d: dout <=  'sd20541; // 893
        'h37e: dout <=  'sd21739; // 894
        'h37f: dout <=  'sd38471; // 895
        'h380: dout <=  'sd48916; // 896
        'h381: dout <= -'sd11964; // 897
        'h382: dout <=  'sd37314; // 898
        'h383: dout <=  'sd19776; // 899
        'h384: dout <=  'sd53096; // 900
        'h385: dout <=  'sd21075; // 901
        'h386: dout <=  'sd4470; // 902
        'h387: dout <=  'sd3768; // 903
        'h388: dout <=  'sd55358; // 904
        'h389: dout <=  'sd4671; // 905
        'h38a: dout <=  'sd41457; // 906
        'h38b: dout <=  'sd43664; // 907
        'h38c: dout <= -'sd52106; // 908
        'h38d: dout <= -'sd42218; // 909
        'h38e: dout <= -'sd2470; // 910
        'h38f: dout <=  'sd48191; // 911
        'h390: dout <= -'sd42905; // 912
        'h391: dout <=  'sd20027; // 913
        'h392: dout <= -'sd44153; // 914
        'h393: dout <=  'sd58554; // 915
        'h394: dout <= -'sd31078; // 916
        'h395: dout <= -'sd52969; // 917
        'h396: dout <= -'sd31584; // 918
        'h397: dout <= -'sd48342; // 919
        'h398: dout <=  'sd39110; // 920
        'h399: dout <=  'sd37507; // 921
        'h39a: dout <=  'sd58592; // 922
        'h39b: dout <=  'sd17699; // 923
        'h39c: dout <=  'sd18499; // 924
        'h39d: dout <=  'sd15135; // 925
        'h39e: dout <=  'sd57992; // 926
        'h39f: dout <=  'sd9907; // 927
        'h3a0: dout <=  'sd56843; // 928
        'h3a1: dout <= -'sd50055; // 929
        'h3a2: dout <= -'sd46675; // 930
        'h3a3: dout <= -'sd21525; // 931
        'h3a4: dout <=  'sd59118; // 932
        'h3a5: dout <= -'sd49877; // 933
        'h3a6: dout <= -'sd16588; // 934
        'h3a7: dout <= -'sd38969; // 935
        'h3a8: dout <=  'sd1944; // 936
        'h3a9: dout <=  'sd1915; // 937
        'h3aa: dout <= -'sd7086; // 938
        'h3ab: dout <=  'sd31354; // 939
        'h3ac: dout <= -'sd549; // 940
        'h3ad: dout <= -'sd59820; // 941
        'h3ae: dout <=  'sd42610; // 942
        'h3af: dout <= -'sd11197; // 943
        'h3b0: dout <=  'sd52756; // 944
        'h3b1: dout <= -'sd55524; // 945
        'h3b2: dout <= -'sd53337; // 946
        'h3b3: dout <=  'sd33124; // 947
        'h3b4: dout <= -'sd42079; // 948
        'h3b5: dout <= -'sd57719; // 949
        'h3b6: dout <= -'sd24687; // 950
        'h3b7: dout <= -'sd2647; // 951
        'h3b8: dout <=  'sd6038; // 952
        'h3b9: dout <=  'sd504; // 953
        'h3ba: dout <=  'sd41704; // 954
        'h3bb: dout <= -'sd23354; // 955
        'h3bc: dout <= -'sd49141; // 956
        'h3bd: dout <= -'sd59631; // 957
        'h3be: dout <= -'sd31497; // 958
        'h3bf: dout <=  'sd40218; // 959
        'h3c0: dout <= -'sd8354; // 960
        'h3c1: dout <= -'sd29281; // 961
        'h3c2: dout <=  'sd14583; // 962
        'h3c3: dout <=  'sd48734; // 963
        'h3c4: dout <=  'sd21263; // 964
        'h3c5: dout <= -'sd21438; // 965
        'h3c6: dout <=  'sd18403; // 966
        'h3c7: dout <= -'sd23133; // 967
        'h3c8: dout <= -'sd39290; // 968
        'h3c9: dout <= -'sd39085; // 969
        'h3ca: dout <= -'sd34815; // 970
        'h3cb: dout <=  'sd20097; // 971
        'h3cc: dout <=  'sd31098; // 972
        'h3cd: dout <=  'sd31528; // 973
        'h3ce: dout <=  'sd117; // 974
        'h3cf: dout <= -'sd11172; // 975
        'h3d0: dout <=  'sd25531; // 976
        'h3d1: dout <=  'sd17355; // 977
        'h3d2: dout <=  'sd58403; // 978
        'h3d3: dout <=  'sd11616; // 979
        'h3d4: dout <= -'sd49454; // 980
        'h3d5: dout <= -'sd52378; // 981
        'h3d6: dout <= -'sd5039; // 982
        'h3d7: dout <= -'sd23282; // 983
        'h3d8: dout <= -'sd10728; // 984
        'h3d9: dout <= -'sd49779; // 985
        'h3da: dout <=  'sd6038; // 986
        'h3db: dout <=  'sd2533; // 987
        'h3dc: dout <= -'sd47874; // 988
        'h3dd: dout <= -'sd30979; // 989
        'h3de: dout <= -'sd48814; // 990
        'h3df: dout <= -'sd3448; // 991
        'h3e0: dout <= -'sd29736; // 992
        'h3e1: dout <= -'sd59987; // 993
        'h3e2: dout <= -'sd40830; // 994
        'h3e3: dout <= -'sd22537; // 995
        'h3e4: dout <= -'sd12246; // 996
        'h3e5: dout <=  'sd38054; // 997
        'h3e6: dout <= -'sd58137; // 998
        'h3e7: dout <=  'sd38899; // 999
        'h3e8: dout <= -'sd57023; // 1000
        'h3e9: dout <=  'sd50644; // 1001
        'h3ea: dout <=  'sd50098; // 1002
        'h3eb: dout <= -'sd49589; // 1003
        'h3ec: dout <= -'sd18163; // 1004
        'h3ed: dout <= -'sd41380; // 1005
        'h3ee: dout <=  'sd54179; // 1006
        'h3ef: dout <=  'sd17865; // 1007
        'h3f0: dout <= -'sd37228; // 1008
        'h3f1: dout <= -'sd4810; // 1009
        'h3f2: dout <= -'sd40371; // 1010
        'h3f3: dout <=  'sd44826; // 1011
        'h3f4: dout <= -'sd11824; // 1012
        'h3f5: dout <=  'sd52382; // 1013
        'h3f6: dout <= -'sd13812; // 1014
        'h3f7: dout <= -'sd20707; // 1015
        'h3f8: dout <= -'sd543; // 1016
        'h3f9: dout <= -'sd48028; // 1017
        'h3fa: dout <= -'sd17207; // 1018
        'h3fb: dout <=  'sd14816; // 1019
        'h3fc: dout <=  'sd12507; // 1020
        'h3fd: dout <=  'sd50418; // 1021
        'h3fe: dout <= -'sd30407; // 1022
        'h3ff: dout <= -'sd22624; // 1023
        'h400: dout <= -'sd46950; // 1024
        'h401: dout <=  'sd37598; // 1025
        'h402: dout <=  'sd41851; // 1026
        'h403: dout <=  'sd43977; // 1027
        'h404: dout <=  'sd21732; // 1028
        'h405: dout <= -'sd35390; // 1029
        'h406: dout <=  'sd1920; // 1030
        'h407: dout <=  'sd59099; // 1031
        'h408: dout <= -'sd7880; // 1032
        'h409: dout <= -'sd45441; // 1033
        'h40a: dout <=  'sd12022; // 1034
        'h40b: dout <=  'sd42820; // 1035
        'h40c: dout <= -'sd28050; // 1036
        'h40d: dout <=  'sd2358; // 1037
        'h40e: dout <= -'sd33251; // 1038
        'h40f: dout <= -'sd45324; // 1039
        'h410: dout <=  'sd25164; // 1040
        'h411: dout <= -'sd47080; // 1041
        'h412: dout <= -'sd54764; // 1042
        'h413: dout <=  'sd18538; // 1043
        'h414: dout <=  'sd37855; // 1044
        'h415: dout <=  'sd43903; // 1045
        'h416: dout <= -'sd22524; // 1046
        'h417: dout <=  'sd46863; // 1047
        'h418: dout <=  'sd37145; // 1048
        'h419: dout <=  'sd17303; // 1049
        'h41a: dout <= -'sd45385; // 1050
        'h41b: dout <=  'sd13443; // 1051
        'h41c: dout <=  'sd58765; // 1052
        'h41d: dout <= -'sd49996; // 1053
        'h41e: dout <= -'sd52863; // 1054
        'h41f: dout <=  'sd57386; // 1055
        'h420: dout <=  'sd34320; // 1056
        'h421: dout <= -'sd55875; // 1057
        'h422: dout <= -'sd28205; // 1058
        'h423: dout <= -'sd17540; // 1059
        'h424: dout <=  'sd43687; // 1060
        'h425: dout <=  'sd29880; // 1061
        'h426: dout <=  'sd34809; // 1062
        'h427: dout <= -'sd30776; // 1063
        'h428: dout <= -'sd59155; // 1064
        'h429: dout <= -'sd30247; // 1065
        'h42a: dout <= -'sd19241; // 1066
        'h42b: dout <=  'sd41163; // 1067
        'h42c: dout <=  'sd34278; // 1068
        'h42d: dout <= -'sd51417; // 1069
        'h42e: dout <=  'sd52071; // 1070
        'h42f: dout <=  'sd44500; // 1071
        'h430: dout <= -'sd42469; // 1072
        'h431: dout <=  'sd47248; // 1073
        'h432: dout <=  'sd58824; // 1074
        'h433: dout <=  'sd57790; // 1075
        'h434: dout <= -'sd36236; // 1076
        'h435: dout <= -'sd5348; // 1077
        'h436: dout <= -'sd3679; // 1078
        'h437: dout <= -'sd20819; // 1079
        'h438: dout <=  'sd45789; // 1080
        'h439: dout <=  'sd55449; // 1081
        'h43a: dout <= -'sd40941; // 1082
        'h43b: dout <=  'sd39921; // 1083
        'h43c: dout <=  'sd14619; // 1084
        'h43d: dout <= -'sd28444; // 1085
        'h43e: dout <= -'sd43084; // 1086
        'h43f: dout <= -'sd9401; // 1087
        'h440: dout <= -'sd60292; // 1088
        'h441: dout <= -'sd34927; // 1089
        'h442: dout <= -'sd14888; // 1090
        'h443: dout <= -'sd18832; // 1091
        'h444: dout <= -'sd47349; // 1092
        'h445: dout <= -'sd1288; // 1093
        'h446: dout <= -'sd11651; // 1094
        'h447: dout <=  'sd59148; // 1095
        'h448: dout <=  'sd49547; // 1096
        'h449: dout <= -'sd20654; // 1097
        'h44a: dout <=  'sd50098; // 1098
        'h44b: dout <=  'sd28427; // 1099
        'h44c: dout <=  'sd47397; // 1100
        'h44d: dout <=  'sd24147; // 1101
        'h44e: dout <=  'sd21788; // 1102
        'h44f: dout <=  'sd47578; // 1103
        'h450: dout <= -'sd22984; // 1104
        'h451: dout <= -'sd1218; // 1105
        'h452: dout <=  'sd54829; // 1106
        'h453: dout <= -'sd49223; // 1107
        'h454: dout <= -'sd15628; // 1108
        'h455: dout <= -'sd38262; // 1109
        'h456: dout <=  'sd2448; // 1110
        'h457: dout <= -'sd50418; // 1111
        'h458: dout <=  'sd45472; // 1112
        'h459: dout <=  'sd1079; // 1113
        'h45a: dout <=  'sd43030; // 1114
        'h45b: dout <= -'sd41534; // 1115
        'h45c: dout <=  'sd49141; // 1116
        'h45d: dout <= -'sd44559; // 1117
        'h45e: dout <=  'sd44519; // 1118
        'h45f: dout <= -'sd45452; // 1119
        'h460: dout <= -'sd47215; // 1120
        'h461: dout <=  'sd35511; // 1121
        'h462: dout <= -'sd23906; // 1122
        'h463: dout <= -'sd12854; // 1123
        'h464: dout <= -'sd6530; // 1124
        'h465: dout <=  'sd20147; // 1125
        'h466: dout <=  'sd9668; // 1126
        'h467: dout <=  'sd45972; // 1127
        'h468: dout <= -'sd36451; // 1128
        'h469: dout <= -'sd58861; // 1129
        'h46a: dout <=  'sd1655; // 1130
        'h46b: dout <= -'sd58453; // 1131
        'h46c: dout <= -'sd48675; // 1132
        'h46d: dout <= -'sd22599; // 1133
        'h46e: dout <=  'sd59268; // 1134
        'h46f: dout <=  'sd56188; // 1135
        'h470: dout <= -'sd57860; // 1136
        'h471: dout <=  'sd8346; // 1137
        'h472: dout <= -'sd15832; // 1138
        'h473: dout <=  'sd37517; // 1139
        'h474: dout <= -'sd55861; // 1140
        'h475: dout <=  'sd40562; // 1141
        'h476: dout <= -'sd37299; // 1142
        'h477: dout <= -'sd43861; // 1143
        'h478: dout <=  'sd13914; // 1144
        'h479: dout <= -'sd11540; // 1145
        'h47a: dout <= -'sd25214; // 1146
        'h47b: dout <= -'sd17269; // 1147
        'h47c: dout <=  'sd8718; // 1148
        'h47d: dout <=  'sd48084; // 1149
        'h47e: dout <=  'sd30229; // 1150
        'h47f: dout <=  'sd51468; // 1151
        'h480: dout <=  'sd19840; // 1152
        'h481: dout <=  'sd52554; // 1153
        'h482: dout <= -'sd38511; // 1154
        'h483: dout <=  'sd964; // 1155
        'h484: dout <= -'sd29344; // 1156
        'h485: dout <= -'sd26787; // 1157
        'h486: dout <=  'sd20967; // 1158
        'h487: dout <= -'sd295; // 1159
        'h488: dout <= -'sd31328; // 1160
        'h489: dout <= -'sd21600; // 1161
        'h48a: dout <= -'sd53393; // 1162
        'h48b: dout <=  'sd46445; // 1163
        'h48c: dout <= -'sd9751; // 1164
        'h48d: dout <=  'sd26555; // 1165
        'h48e: dout <= -'sd49533; // 1166
        'h48f: dout <= -'sd39385; // 1167
        'h490: dout <= -'sd22295; // 1168
        'h491: dout <= -'sd46056; // 1169
        'h492: dout <=  'sd12729; // 1170
        'h493: dout <=  'sd23404; // 1171
        'h494: dout <= -'sd5422; // 1172
        'h495: dout <= -'sd10013; // 1173
        'h496: dout <= -'sd875; // 1174
        'h497: dout <= -'sd54318; // 1175
        'h498: dout <= -'sd20407; // 1176
        'h499: dout <= -'sd58043; // 1177
        'h49a: dout <=  'sd29900; // 1178
        'h49b: dout <=  'sd27009; // 1179
        'h49c: dout <= -'sd16842; // 1180
        'h49d: dout <=  'sd16217; // 1181
        'h49e: dout <= -'sd39988; // 1182
        'h49f: dout <= -'sd14824; // 1183
        'h4a0: dout <= -'sd51633; // 1184
        'h4a1: dout <= -'sd32884; // 1185
        'h4a2: dout <= -'sd12919; // 1186
        'h4a3: dout <= -'sd16424; // 1187
        'h4a4: dout <= -'sd43221; // 1188
        'h4a5: dout <= -'sd59761; // 1189
        'h4a6: dout <= -'sd16387; // 1190
        'h4a7: dout <=  'sd59155; // 1191
        'h4a8: dout <= -'sd53762; // 1192
        'h4a9: dout <=  'sd58579; // 1193
        'h4aa: dout <= -'sd32201; // 1194
        'h4ab: dout <=  'sd29441; // 1195
        'h4ac: dout <= -'sd8731; // 1196
        'h4ad: dout <=  'sd1078; // 1197
        'h4ae: dout <=  'sd51431; // 1198
        'h4af: dout <=  'sd5732; // 1199
        'h4b0: dout <=  'sd23182; // 1200
        'h4b1: dout <= -'sd36157; // 1201
        'h4b2: dout <=  'sd3038; // 1202
        'h4b3: dout <= -'sd24548; // 1203
        'h4b4: dout <= -'sd52217; // 1204
        'h4b5: dout <= -'sd9517; // 1205
        'h4b6: dout <= -'sd56347; // 1206
        'h4b7: dout <= -'sd33803; // 1207
        'h4b8: dout <= -'sd59195; // 1208
        'h4b9: dout <=  'sd55005; // 1209
        'h4ba: dout <= -'sd55185; // 1210
        'h4bb: dout <= -'sd44741; // 1211
        'h4bc: dout <= -'sd37177; // 1212
        'h4bd: dout <=  'sd32328; // 1213
        'h4be: dout <=  'sd9185; // 1214
        'h4bf: dout <=  'sd25271; // 1215
        'h4c0: dout <= -'sd8660; // 1216
        'h4c1: dout <= -'sd6951; // 1217
        'h4c2: dout <= -'sd18543; // 1218
        'h4c3: dout <=  'sd20288; // 1219
        'h4c4: dout <=  'sd35128; // 1220
        'h4c5: dout <=  'sd51823; // 1221
        'h4c6: dout <=  'sd5396; // 1222
        'h4c7: dout <=  'sd41633; // 1223
        'h4c8: dout <=  'sd713; // 1224
        'h4c9: dout <= -'sd51012; // 1225
        'h4ca: dout <=  'sd51881; // 1226
        'h4cb: dout <= -'sd16491; // 1227
        'h4cc: dout <= -'sd56651; // 1228
        'h4cd: dout <=  'sd37356; // 1229
        'h4ce: dout <=  'sd4704; // 1230
        'h4cf: dout <=  'sd45760; // 1231
        'h4d0: dout <=  'sd16490; // 1232
        'h4d1: dout <=  'sd49918; // 1233
        'h4d2: dout <=  'sd26425; // 1234
        'h4d3: dout <=  'sd15284; // 1235
        'h4d4: dout <=  'sd38569; // 1236
        'h4d5: dout <= -'sd51879; // 1237
        'h4d6: dout <= -'sd38708; // 1238
        'h4d7: dout <= -'sd15454; // 1239
        'h4d8: dout <=  'sd41458; // 1240
        'h4d9: dout <=  'sd44746; // 1241
        'h4da: dout <=  'sd44325; // 1242
        'h4db: dout <=  'sd3237; // 1243
        'h4dc: dout <= -'sd30918; // 1244
        'h4dd: dout <= -'sd3862; // 1245
        'h4de: dout <= -'sd17988; // 1246
        'h4df: dout <= -'sd12644; // 1247
        'h4e0: dout <= -'sd30018; // 1248
        'h4e1: dout <= -'sd17814; // 1249
        'h4e2: dout <=  'sd5881; // 1250
        'h4e3: dout <= -'sd10256; // 1251
        'h4e4: dout <=  'sd44902; // 1252
        'h4e5: dout <= -'sd5665; // 1253
        'h4e6: dout <=  'sd4623; // 1254
        'h4e7: dout <= -'sd49192; // 1255
        'h4e8: dout <= -'sd20660; // 1256
        'h4e9: dout <= -'sd42507; // 1257
        'h4ea: dout <= -'sd28986; // 1258
        'h4eb: dout <= -'sd23593; // 1259
        'h4ec: dout <=  'sd5990; // 1260
        'h4ed: dout <=  'sd3904; // 1261
        'h4ee: dout <=  'sd20284; // 1262
        'h4ef: dout <= -'sd59989; // 1263
        'h4f0: dout <= -'sd55256; // 1264
        'h4f1: dout <=  'sd14370; // 1265
        'h4f2: dout <= -'sd51383; // 1266
        'h4f3: dout <= -'sd19597; // 1267
        'h4f4: dout <=  'sd39192; // 1268
        'h4f5: dout <=  'sd20936; // 1269
        'h4f6: dout <=  'sd28931; // 1270
        'h4f7: dout <= -'sd36680; // 1271
        'h4f8: dout <= -'sd58618; // 1272
        'h4f9: dout <=  'sd42622; // 1273
        'h4fa: dout <= -'sd28657; // 1274
        'h4fb: dout <= -'sd16070; // 1275
        'h4fc: dout <= -'sd24751; // 1276
        'h4fd: dout <= -'sd24858; // 1277
        'h4fe: dout <= -'sd18645; // 1278
        'h4ff: dout <=  'sd10247; // 1279
        'h500: dout <=  'sd4345; // 1280
        'h501: dout <=  'sd18992; // 1281
        'h502: dout <= -'sd32833; // 1282
        'h503: dout <= -'sd35573; // 1283
        'h504: dout <=  'sd22947; // 1284
        'h505: dout <=  'sd54597; // 1285
        'h506: dout <=  'sd34887; // 1286
        'h507: dout <= -'sd41669; // 1287
        'h508: dout <= -'sd22216; // 1288
        'h509: dout <=  'sd8704; // 1289
        'h50a: dout <= -'sd20024; // 1290
        'h50b: dout <= -'sd35290; // 1291
        'h50c: dout <=  'sd23673; // 1292
        'h50d: dout <=  'sd38374; // 1293
        'h50e: dout <=  'sd51379; // 1294
        'h50f: dout <= -'sd26445; // 1295
        'h510: dout <= -'sd30386; // 1296
        'h511: dout <= -'sd15005; // 1297
        'h512: dout <=  'sd47730; // 1298
        'h513: dout <= -'sd59636; // 1299
        'h514: dout <=  'sd19664; // 1300
        'h515: dout <=  'sd34636; // 1301
        'h516: dout <= -'sd23164; // 1302
        'h517: dout <=  'sd34890; // 1303
        'h518: dout <=  'sd15207; // 1304
        'h519: dout <=  'sd25374; // 1305
        'h51a: dout <=  'sd12532; // 1306
        'h51b: dout <= -'sd32675; // 1307
        'h51c: dout <=  'sd45909; // 1308
        'h51d: dout <=  'sd23928; // 1309
        'h51e: dout <= -'sd47171; // 1310
        'h51f: dout <=  'sd36751; // 1311
        'h520: dout <= -'sd11925; // 1312
        'h521: dout <= -'sd396; // 1313
        'h522: dout <=  'sd44001; // 1314
        'h523: dout <= -'sd36692; // 1315
        'h524: dout <=  'sd50271; // 1316
        'h525: dout <= -'sd57489; // 1317
        'h526: dout <= -'sd37896; // 1318
        'h527: dout <=  'sd45585; // 1319
        'h528: dout <= -'sd49332; // 1320
        'h529: dout <= -'sd30311; // 1321
        'h52a: dout <=  'sd28867; // 1322
        'h52b: dout <= -'sd31681; // 1323
        'h52c: dout <= -'sd41606; // 1324
        'h52d: dout <= -'sd33476; // 1325
        'h52e: dout <=  'sd57727; // 1326
        'h52f: dout <= -'sd39928; // 1327
        'h530: dout <=  'sd19007; // 1328
        'h531: dout <= -'sd50946; // 1329
        'h532: dout <=  'sd50838; // 1330
        'h533: dout <=  'sd8742; // 1331
        'h534: dout <= -'sd6804; // 1332
        'h535: dout <=  'sd59474; // 1333
        'h536: dout <= -'sd16010; // 1334
        'h537: dout <= -'sd27027; // 1335
        'h538: dout <=  'sd33034; // 1336
        'h539: dout <=  'sd4986; // 1337
        'h53a: dout <=  'sd59304; // 1338
        'h53b: dout <=  'sd12908; // 1339
        'h53c: dout <= -'sd45673; // 1340
        'h53d: dout <= -'sd34883; // 1341
        'h53e: dout <=  'sd23299; // 1342
        'h53f: dout <= -'sd51236; // 1343
        'h540: dout <=  'sd56952; // 1344
        'h541: dout <= -'sd429; // 1345
        'h542: dout <= -'sd32058; // 1346
        'h543: dout <=  'sd28862; // 1347
        'h544: dout <=  'sd3203; // 1348
        'h545: dout <= -'sd28793; // 1349
        'h546: dout <= -'sd5630; // 1350
        'h547: dout <= -'sd53305; // 1351
        'h548: dout <=  'sd48159; // 1352
        'h549: dout <= -'sd1153; // 1353
        'h54a: dout <= -'sd43896; // 1354
        'h54b: dout <= -'sd46399; // 1355
        'h54c: dout <= -'sd36848; // 1356
        'h54d: dout <= -'sd7475; // 1357
        'h54e: dout <=  'sd35959; // 1358
        'h54f: dout <= -'sd42292; // 1359
        'h550: dout <= -'sd57838; // 1360
        'h551: dout <= -'sd1620; // 1361
        'h552: dout <=  'sd2589; // 1362
        'h553: dout <=  'sd58512; // 1363
        'h554: dout <=  'sd25515; // 1364
        'h555: dout <=  'sd43525; // 1365
        'h556: dout <= -'sd54524; // 1366
        'h557: dout <= -'sd41676; // 1367
        'h558: dout <=  'sd39412; // 1368
        'h559: dout <= -'sd47472; // 1369
        'h55a: dout <=  'sd38909; // 1370
        'h55b: dout <= -'sd20840; // 1371
        'h55c: dout <=  'sd7841; // 1372
        'h55d: dout <= -'sd42088; // 1373
        'h55e: dout <=  'sd6793; // 1374
        'h55f: dout <= -'sd14290; // 1375
        'h560: dout <= -'sd51496; // 1376
        'h561: dout <=  'sd43226; // 1377
        'h562: dout <=  'sd26292; // 1378
        'h563: dout <=  'sd19317; // 1379
        'h564: dout <=  'sd33586; // 1380
        'h565: dout <= -'sd16187; // 1381
        'h566: dout <= -'sd10575; // 1382
        'h567: dout <=  'sd48328; // 1383
        'h568: dout <= -'sd32444; // 1384
        'h569: dout <=  'sd22700; // 1385
        'h56a: dout <= -'sd5888; // 1386
        'h56b: dout <=  'sd19950; // 1387
        'h56c: dout <= -'sd51787; // 1388
        'h56d: dout <= -'sd19482; // 1389
        'h56e: dout <=  'sd9947; // 1390
        'h56f: dout <= -'sd57380; // 1391
        'h570: dout <=  'sd2896; // 1392
        'h571: dout <= -'sd4805; // 1393
        'h572: dout <= -'sd630; // 1394
        'h573: dout <=  'sd31377; // 1395
        'h574: dout <=  'sd43266; // 1396
        'h575: dout <=  'sd18136; // 1397
        'h576: dout <= -'sd58345; // 1398
        'h577: dout <=  'sd8461; // 1399
        'h578: dout <= -'sd27130; // 1400
        'h579: dout <= -'sd45723; // 1401
        'h57a: dout <= -'sd44784; // 1402
        'h57b: dout <= -'sd32089; // 1403
        'h57c: dout <=  'sd58426; // 1404
        'h57d: dout <= -'sd19289; // 1405
        'h57e: dout <= -'sd117; // 1406
        'h57f: dout <=  'sd44291; // 1407
        'h580: dout <=  'sd14653; // 1408
        'h581: dout <=  'sd50588; // 1409
        'h582: dout <=  'sd4404; // 1410
        'h583: dout <=  'sd9384; // 1411
        'h584: dout <=  'sd32410; // 1412
        'h585: dout <=  'sd49864; // 1413
        'h586: dout <=  'sd18384; // 1414
        'h587: dout <= -'sd37941; // 1415
        'h588: dout <=  'sd35645; // 1416
        'h589: dout <=  'sd58832; // 1417
        'h58a: dout <=  'sd10316; // 1418
        'h58b: dout <= -'sd36621; // 1419
        'h58c: dout <= -'sd7917; // 1420
        'h58d: dout <=  'sd34575; // 1421
        'h58e: dout <= -'sd18234; // 1422
        'h58f: dout <= -'sd24145; // 1423
        'h590: dout <=  'sd34979; // 1424
        'h591: dout <=  'sd11883; // 1425
        'h592: dout <=  'sd49745; // 1426
        'h593: dout <= -'sd13693; // 1427
        'h594: dout <=  'sd10802; // 1428
        'h595: dout <= -'sd5926; // 1429
        'h596: dout <= -'sd12845; // 1430
        'h597: dout <= -'sd6086; // 1431
        'h598: dout <= -'sd6463; // 1432
        'h599: dout <= -'sd28787; // 1433
        'h59a: dout <=  'sd53609; // 1434
        'h59b: dout <=  'sd45240; // 1435
        'h59c: dout <=  'sd14024; // 1436
        'h59d: dout <= -'sd15784; // 1437
        'h59e: dout <= -'sd49777; // 1438
        'h59f: dout <=  'sd51994; // 1439
        'h5a0: dout <= -'sd26262; // 1440
        'h5a1: dout <=  'sd19693; // 1441
        'h5a2: dout <= -'sd59887; // 1442
        'h5a3: dout <= -'sd10604; // 1443
        'h5a4: dout <=  'sd52173; // 1444
        'h5a5: dout <= -'sd32969; // 1445
        'h5a6: dout <=  'sd24911; // 1446
        'h5a7: dout <= -'sd38660; // 1447
        'h5a8: dout <=  'sd25063; // 1448
        'h5a9: dout <=  'sd7391; // 1449
        'h5aa: dout <=  'sd16425; // 1450
        'h5ab: dout <=  'sd21630; // 1451
        'h5ac: dout <= -'sd10542; // 1452
        'h5ad: dout <= -'sd19527; // 1453
        'h5ae: dout <= -'sd44751; // 1454
        'h5af: dout <=  'sd7335; // 1455
        'h5b0: dout <=  'sd16531; // 1456
        'h5b1: dout <=  'sd9534; // 1457
        'h5b2: dout <= -'sd35660; // 1458
        'h5b3: dout <=  'sd9208; // 1459
        'h5b4: dout <=  'sd45288; // 1460
        'h5b5: dout <= -'sd6560; // 1461
        'h5b6: dout <= -'sd49931; // 1462
        'h5b7: dout <= -'sd60318; // 1463
        'h5b8: dout <=  'sd33630; // 1464
        'h5b9: dout <=  'sd46159; // 1465
        'h5ba: dout <=  'sd36222; // 1466
        'h5bb: dout <=  'sd45534; // 1467
        'h5bc: dout <=  'sd15231; // 1468
        'h5bd: dout <= -'sd29884; // 1469
        'h5be: dout <=  'sd6246; // 1470
        'h5bf: dout <=  'sd16349; // 1471
        'h5c0: dout <= -'sd51289; // 1472
        'h5c1: dout <= -'sd4912; // 1473
        'h5c2: dout <=  'sd29094; // 1474
        'h5c3: dout <= -'sd34350; // 1475
        'h5c4: dout <= -'sd49634; // 1476
        'h5c5: dout <=  'sd41701; // 1477
        'h5c6: dout <=  'sd55944; // 1478
        'h5c7: dout <=  'sd25896; // 1479
        'h5c8: dout <= -'sd56938; // 1480
        'h5c9: dout <= -'sd52885; // 1481
        'h5ca: dout <=  'sd12857; // 1482
        'h5cb: dout <=  'sd30065; // 1483
        'h5cc: dout <= -'sd54845; // 1484
        'h5cd: dout <=  'sd29611; // 1485
        'h5ce: dout <=  'sd34354; // 1486
        'h5cf: dout <= -'sd3051; // 1487
        'h5d0: dout <= -'sd30712; // 1488
        'h5d1: dout <=  'sd47683; // 1489
        'h5d2: dout <=  'sd48782; // 1490
        'h5d3: dout <=  'sd32349; // 1491
        'h5d4: dout <=  'sd31088; // 1492
        'h5d5: dout <= -'sd4240; // 1493
        'h5d6: dout <= -'sd50816; // 1494
        'h5d7: dout <= -'sd17818; // 1495
        'h5d8: dout <= -'sd20198; // 1496
        'h5d9: dout <=  'sd18982; // 1497
        'h5da: dout <= -'sd48358; // 1498
        'h5db: dout <= -'sd990; // 1499
        'h5dc: dout <=  'sd58239; // 1500
        'h5dd: dout <= -'sd40299; // 1501
        'h5de: dout <=  'sd35893; // 1502
        'h5df: dout <= -'sd34298; // 1503
        'h5e0: dout <=  'sd14338; // 1504
        'h5e1: dout <=  'sd3467; // 1505
        'h5e2: dout <= -'sd17390; // 1506
        'h5e3: dout <=  'sd1934; // 1507
        'h5e4: dout <=  'sd34360; // 1508
        'h5e5: dout <= -'sd24540; // 1509
        'h5e6: dout <= -'sd23026; // 1510
        'h5e7: dout <= -'sd13318; // 1511
        'h5e8: dout <=  'sd31689; // 1512
        'h5e9: dout <= -'sd22941; // 1513
        'h5ea: dout <= -'sd38186; // 1514
        'h5eb: dout <=  'sd55964; // 1515
        'h5ec: dout <=  'sd26726; // 1516
        'h5ed: dout <= -'sd3507; // 1517
        'h5ee: dout <= -'sd8047; // 1518
        'h5ef: dout <=  'sd53946; // 1519
        'h5f0: dout <= -'sd5636; // 1520
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

