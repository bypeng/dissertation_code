module mod4621Svec33 (
    input       [32:0] z_in,
    output      [11:0] p0,
    output reg  [11:0] p1,
    output reg  [11:0] p2,
    output reg  [11:0] p3,
    output reg  [11:0] n0,
    output reg  [12:0] n1
) ;

    assign p0 = z_in[11:0];

    always @ (*) begin
        case({ z_in[27], z_in[16], z_in[15] })
            3'h0: p1 = 12'd0;
            3'h1: p1 = 12'd421;
            3'h2: p1 = 12'd842;
            3'h3: p1 = 12'd1263;
            3'h4: p1 = 12'd783;
            3'h5: p1 = 12'd1204;
            3'h6: p1 = 12'd1625;
            3'h7: p1 = 12'd2046;
        endcase
    end

    always @ (*) begin
        case({ z_in[31], z_in[30], z_in[28], z_in[23], z_in[18], z_in[17] })
            6'h00: p2 = 12'd0;
            6'h01: p2 = 12'd1684;
            6'h02: p2 = 12'd3368;
            6'h03: p2 = 12'd431;
            6'h04: p2 = 12'd1493;
            6'h05: p2 = 12'd3177;
            6'h06: p2 = 12'd240;
            6'h07: p2 = 12'd1924;
            6'h08: p2 = 12'd1566;
            6'h09: p2 = 12'd3250;
            6'h0a: p2 = 12'd313;
            6'h0b: p2 = 12'd1997;
            6'h0c: p2 = 12'd3059;
            6'h0d: p2 = 12'd122;
            6'h0e: p2 = 12'd1806;
            6'h0f: p2 = 12'd3490;
            6'h10: p2 = 12'd1643;
            6'h11: p2 = 12'd3327;
            6'h12: p2 = 12'd390;
            6'h13: p2 = 12'd2074;
            6'h14: p2 = 12'd3136;
            6'h15: p2 = 12'd199;
            6'h16: p2 = 12'd1883;
            6'h17: p2 = 12'd3567;
            6'h18: p2 = 12'd3209;
            6'h19: p2 = 12'd272;
            6'h1a: p2 = 12'd1956;
            6'h1b: p2 = 12'd3640;
            6'h1c: p2 = 12'd81;
            6'h1d: p2 = 12'd1765;
            6'h1e: p2 = 12'd3449;
            6'h1f: p2 = 12'd512;
            6'h20: p2 = 12'd3286;
            6'h21: p2 = 12'd349;
            6'h22: p2 = 12'd2033;
            6'h23: p2 = 12'd3717;
            6'h24: p2 = 12'd158;
            6'h25: p2 = 12'd1842;
            6'h26: p2 = 12'd3526;
            6'h27: p2 = 12'd589;
            6'h28: p2 = 12'd231;
            6'h29: p2 = 12'd1915;
            6'h2a: p2 = 12'd3599;
            6'h2b: p2 = 12'd662;
            6'h2c: p2 = 12'd1724;
            6'h2d: p2 = 12'd3408;
            6'h2e: p2 = 12'd471;
            6'h2f: p2 = 12'd2155;
            6'h30: p2 = 12'd308;
            6'h31: p2 = 12'd1992;
            6'h32: p2 = 12'd3676;
            6'h33: p2 = 12'd739;
            6'h34: p2 = 12'd1801;
            6'h35: p2 = 12'd3485;
            6'h36: p2 = 12'd548;
            6'h37: p2 = 12'd2232;
            6'h38: p2 = 12'd1874;
            6'h39: p2 = 12'd3558;
            6'h3a: p2 = 12'd621;
            6'h3b: p2 = 12'd2305;
            6'h3c: p2 = 12'd3367;
            6'h3d: p2 = 12'd430;
            6'h3e: p2 = 12'd2114;
            6'h3f: p2 = 12'd3798;
        endcase
    end

    always @ (*) begin
        case({ z_in[32], z_in[19], z_in[14] })
            3'h0: p3 = 12'd0;
            3'h1: p3 = 12'd2521;
            3'h2: p3 = 12'd2115;
            3'h3: p3 = 12'd15;
            3'h4: p3 = 12'd2670;
            3'h5: p3 = 12'd570;
            3'h6: p3 = 12'd164;
            3'h7: p3 = 12'd2685;
        endcase
    end

    always @ (*) begin
        case({ z_in[21], z_in[13], z_in[12] })
            3'h0: n0 = 12'd0;
            3'h1: n0 = 12'd525;
            3'h2: n0 = 12'd1050;
            3'h3: n0 = 12'd1575;
            3'h4: n0 = 12'd782;
            3'h5: n0 = 12'd1307;
            3'h6: n0 = 12'd1832;
            3'h7: n0 = 12'd2357;
        endcase
    end

    always @ (*) begin
        case({ z_in[29], z_in[26], z_in[25], z_in[24], z_in[22], z_in[20] })
            6'h00: n1 = 13'd0;
            6'h01: n1 = 13'd391;
            6'h02: n1 = 13'd1564;
            6'h03: n1 = 13'd1955;
            6'h04: n1 = 13'd1635;
            6'h05: n1 = 13'd2026;
            6'h06: n1 = 13'd3199;
            6'h07: n1 = 13'd3590;
            6'h08: n1 = 13'd3270;
            6'h09: n1 = 13'd3661;
            6'h0a: n1 = 13'd213;
            6'h0b: n1 = 13'd604;
            6'h0c: n1 = 13'd284;
            6'h0d: n1 = 13'd675;
            6'h0e: n1 = 13'd1848;
            6'h0f: n1 = 13'd2239;
            6'h10: n1 = 13'd1919;
            6'h11: n1 = 13'd2310;
            6'h12: n1 = 13'd3483;
            6'h13: n1 = 13'd3874;
            6'h14: n1 = 13'd3554;
            6'h15: n1 = 13'd3945;
            6'h16: n1 = 13'd497;
            6'h17: n1 = 13'd888;
            6'h18: n1 = 13'd568;
            6'h19: n1 = 13'd959;
            6'h1a: n1 = 13'd2132;
            6'h1b: n1 = 13'd2523;
            6'h1c: n1 = 13'd2203;
            6'h1d: n1 = 13'd2594;
            6'h1e: n1 = 13'd3767;
            6'h1f: n1 = 13'd4158;
            6'h20: n1 = 13'd1489;
            6'h21: n1 = 13'd1880;
            6'h22: n1 = 13'd3053;
            6'h23: n1 = 13'd3444;
            6'h24: n1 = 13'd3124;
            6'h25: n1 = 13'd3515;
            6'h26: n1 = 13'd67;
            6'h27: n1 = 13'd458;
            6'h28: n1 = 13'd138;
            6'h29: n1 = 13'd529;
            6'h2a: n1 = 13'd1702;
            6'h2b: n1 = 13'd2093;
            6'h2c: n1 = 13'd1773;
            6'h2d: n1 = 13'd2164;
            6'h2e: n1 = 13'd3337;
            6'h2f: n1 = 13'd3728;
            6'h30: n1 = 13'd3408;
            6'h31: n1 = 13'd3799;
            6'h32: n1 = 13'd351;
            6'h33: n1 = 13'd742;
            6'h34: n1 = 13'd422;
            6'h35: n1 = 13'd813;
            6'h36: n1 = 13'd1986;
            6'h37: n1 = 13'd2377;
            6'h38: n1 = 13'd2057;
            6'h39: n1 = 13'd2448;
            6'h3a: n1 = 13'd3621;
            6'h3b: n1 = 13'd4012;
            6'h3c: n1 = 13'd3692;
            6'h3d: n1 = 13'd4083;
            6'h3e: n1 = 13'd635;
            6'h3f: n1 = 13'd1026;
        endcase
    end

endmodule
