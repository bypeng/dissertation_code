module mem_ref ( clk, in_addr, in_data, out_addr, out_data_ref ) ;

  localparam DS_CNT = 'd1;
  localparam DS_DEPTH = 'd0;
  localparam B_LEN = 'd1317;
  localparam B_DEPTH = 'd11;
  localparam R_LEN = 'd953;
  localparam R_DEPTH = 'd10;

  input              clk;
  input      [10: 0] in_addr;
  output reg [ 7: 0] in_data;
  input      [ 9: 0] out_addr;
  output reg [13: 0] out_data_ref;

  always @ ( posedge clk ) begin
    case(in_addr)
      11'd0    : in_data <= 8'h6a;
      11'd1    : in_data <= 8'hc8;
      11'd2    : in_data <= 8'hfa;
      11'd3    : in_data <= 8'hd2;
      11'd4    : in_data <= 8'hc3;
      11'd5    : in_data <= 8'h21;
      11'd6    : in_data <= 8'h1a;
      11'd7    : in_data <= 8'h24;
      11'd8    : in_data <= 8'heb;
      11'd9    : in_data <= 8'hf1;
      11'd10   : in_data <= 8'hbd;
      11'd11   : in_data <= 8'h34;
      11'd12   : in_data <= 8'hf4;
      11'd13   : in_data <= 8'h26;
      11'd14   : in_data <= 8'h08;
      11'd15   : in_data <= 8'hf2;
      11'd16   : in_data <= 8'h76;
      11'd17   : in_data <= 8'h27;
      11'd18   : in_data <= 8'h42;
      11'd19   : in_data <= 8'heb;
      11'd20   : in_data <= 8'h7f;
      11'd21   : in_data <= 8'h0b;
      11'd22   : in_data <= 8'h29;
      11'd23   : in_data <= 8'hca;
      11'd24   : in_data <= 8'he6;
      11'd25   : in_data <= 8'hae;
      11'd26   : in_data <= 8'hfc;
      11'd27   : in_data <= 8'h11;
      11'd28   : in_data <= 8'h78;
      11'd29   : in_data <= 8'hdf;
      11'd30   : in_data <= 8'h30;
      11'd31   : in_data <= 8'h90;
      11'd32   : in_data <= 8'h6d;
      11'd33   : in_data <= 8'h75;
      11'd34   : in_data <= 8'hb7;
      11'd35   : in_data <= 8'ha7;
      11'd36   : in_data <= 8'h3b;
      11'd37   : in_data <= 8'h1f;
      11'd38   : in_data <= 8'h33;
      11'd39   : in_data <= 8'h44;
      11'd40   : in_data <= 8'he5;
      11'd41   : in_data <= 8'h6d;
      11'd42   : in_data <= 8'hb9;
      11'd43   : in_data <= 8'hf8;
      11'd44   : in_data <= 8'h55;
      11'd45   : in_data <= 8'h74;
      11'd46   : in_data <= 8'h89;
      11'd47   : in_data <= 8'ha5;
      11'd48   : in_data <= 8'haf;
      11'd49   : in_data <= 8'h60;
      11'd50   : in_data <= 8'had;
      11'd51   : in_data <= 8'h91;
      11'd52   : in_data <= 8'h10;
      11'd53   : in_data <= 8'h52;
      11'd54   : in_data <= 8'h43;
      11'd55   : in_data <= 8'h2f;
      11'd56   : in_data <= 8'he9;
      11'd57   : in_data <= 8'h31;
      11'd58   : in_data <= 8'h56;
      11'd59   : in_data <= 8'h8d;
      11'd60   : in_data <= 8'h3d;
      11'd61   : in_data <= 8'hd0;
      11'd62   : in_data <= 8'hd9;
      11'd63   : in_data <= 8'h18;
      11'd64   : in_data <= 8'h4a;
      11'd65   : in_data <= 8'hf9;
      11'd66   : in_data <= 8'h45;
      11'd67   : in_data <= 8'h3b;
      11'd68   : in_data <= 8'hb3;
      11'd69   : in_data <= 8'h44;
      11'd70   : in_data <= 8'h54;
      11'd71   : in_data <= 8'h8f;
      11'd72   : in_data <= 8'hbf;
      11'd73   : in_data <= 8'h76;
      11'd74   : in_data <= 8'hd8;
      11'd75   : in_data <= 8'h10;
      11'd76   : in_data <= 8'hb3;
      11'd77   : in_data <= 8'h09;
      11'd78   : in_data <= 8'h32;
      11'd79   : in_data <= 8'hfd;
      11'd80   : in_data <= 8'ha7;
      11'd81   : in_data <= 8'h68;
      11'd82   : in_data <= 8'hb4;
      11'd83   : in_data <= 8'h6d;
      11'd84   : in_data <= 8'he9;
      11'd85   : in_data <= 8'h71;
      11'd86   : in_data <= 8'hb4;
      11'd87   : in_data <= 8'hd4;
      11'd88   : in_data <= 8'h35;
      11'd89   : in_data <= 8'h06;
      11'd90   : in_data <= 8'h45;
      11'd91   : in_data <= 8'h62;
      11'd92   : in_data <= 8'hfb;
      11'd93   : in_data <= 8'he2;
      11'd94   : in_data <= 8'h52;
      11'd95   : in_data <= 8'h50;
      11'd96   : in_data <= 8'h79;
      11'd97   : in_data <= 8'hd5;
      11'd98   : in_data <= 8'hf9;
      11'd99   : in_data <= 8'hbc;
      11'd100  : in_data <= 8'hef;
      11'd101  : in_data <= 8'h57;
      11'd102  : in_data <= 8'h21;
      11'd103  : in_data <= 8'h20;
      11'd104  : in_data <= 8'hef;
      11'd105  : in_data <= 8'h4e;
      11'd106  : in_data <= 8'h0c;
      11'd107  : in_data <= 8'h6d;
      11'd108  : in_data <= 8'h84;
      11'd109  : in_data <= 8'hb9;
      11'd110  : in_data <= 8'h25;
      11'd111  : in_data <= 8'h5f;
      11'd112  : in_data <= 8'hf6;
      11'd113  : in_data <= 8'h16;
      11'd114  : in_data <= 8'hbc;
      11'd115  : in_data <= 8'h05;
      11'd116  : in_data <= 8'hcc;
      11'd117  : in_data <= 8'h25;
      11'd118  : in_data <= 8'he0;
      11'd119  : in_data <= 8'h45;
      11'd120  : in_data <= 8'hac;
      11'd121  : in_data <= 8'h25;
      11'd122  : in_data <= 8'hcf;
      11'd123  : in_data <= 8'hb9;
      11'd124  : in_data <= 8'hca;
      11'd125  : in_data <= 8'h3f;
      11'd126  : in_data <= 8'hd3;
      11'd127  : in_data <= 8'h3a;
      11'd128  : in_data <= 8'h4f;
      11'd129  : in_data <= 8'h1d;
      11'd130  : in_data <= 8'h81;
      11'd131  : in_data <= 8'hb2;
      11'd132  : in_data <= 8'h2b;
      11'd133  : in_data <= 8'h1c;
      11'd134  : in_data <= 8'h9d;
      11'd135  : in_data <= 8'h21;
      11'd136  : in_data <= 8'hf7;
      11'd137  : in_data <= 8'hd0;
      11'd138  : in_data <= 8'h6f;
      11'd139  : in_data <= 8'h9b;
      11'd140  : in_data <= 8'h0d;
      11'd141  : in_data <= 8'h9b;
      11'd142  : in_data <= 8'h50;
      11'd143  : in_data <= 8'h12;
      11'd144  : in_data <= 8'h6e;
      11'd145  : in_data <= 8'he7;
      11'd146  : in_data <= 8'h5f;
      11'd147  : in_data <= 8'h45;
      11'd148  : in_data <= 8'h55;
      11'd149  : in_data <= 8'h6a;
      11'd150  : in_data <= 8'ha6;
      11'd151  : in_data <= 8'hf3;
      11'd152  : in_data <= 8'hb3;
      11'd153  : in_data <= 8'h97;
      11'd154  : in_data <= 8'h7b;
      11'd155  : in_data <= 8'hde;
      11'd156  : in_data <= 8'hd6;
      11'd157  : in_data <= 8'h94;
      11'd158  : in_data <= 8'hc2;
      11'd159  : in_data <= 8'h39;
      11'd160  : in_data <= 8'h67;
      11'd161  : in_data <= 8'h4b;
      11'd162  : in_data <= 8'h0f;
      11'd163  : in_data <= 8'h92;
      11'd164  : in_data <= 8'h4b;
      11'd165  : in_data <= 8'h87;
      11'd166  : in_data <= 8'hd9;
      11'd167  : in_data <= 8'h89;
      11'd168  : in_data <= 8'hf6;
      11'd169  : in_data <= 8'h73;
      11'd170  : in_data <= 8'h24;
      11'd171  : in_data <= 8'h95;
      11'd172  : in_data <= 8'h0b;
      11'd173  : in_data <= 8'hd8;
      11'd174  : in_data <= 8'hfb;
      11'd175  : in_data <= 8'h38;
      11'd176  : in_data <= 8'hf0;
      11'd177  : in_data <= 8'h54;
      11'd178  : in_data <= 8'h65;
      11'd179  : in_data <= 8'hce;
      11'd180  : in_data <= 8'hb7;
      11'd181  : in_data <= 8'he4;
      11'd182  : in_data <= 8'hf7;
      11'd183  : in_data <= 8'hd7;
      11'd184  : in_data <= 8'he1;
      11'd185  : in_data <= 8'h3d;
      11'd186  : in_data <= 8'he5;
      11'd187  : in_data <= 8'h16;
      11'd188  : in_data <= 8'hcf;
      11'd189  : in_data <= 8'h71;
      11'd190  : in_data <= 8'h1c;
      11'd191  : in_data <= 8'h58;
      11'd192  : in_data <= 8'h24;
      11'd193  : in_data <= 8'ha0;
      11'd194  : in_data <= 8'h2a;
      11'd195  : in_data <= 8'h56;
      11'd196  : in_data <= 8'hc7;
      11'd197  : in_data <= 8'h1f;
      11'd198  : in_data <= 8'h55;
      11'd199  : in_data <= 8'h58;
      11'd200  : in_data <= 8'h2e;
      11'd201  : in_data <= 8'ha0;
      11'd202  : in_data <= 8'h55;
      11'd203  : in_data <= 8'h8e;
      11'd204  : in_data <= 8'h9b;
      11'd205  : in_data <= 8'h81;
      11'd206  : in_data <= 8'hef;
      11'd207  : in_data <= 8'h08;
      11'd208  : in_data <= 8'h5a;
      11'd209  : in_data <= 8'h7f;
      11'd210  : in_data <= 8'h7e;
      11'd211  : in_data <= 8'h29;
      11'd212  : in_data <= 8'h3e;
      11'd213  : in_data <= 8'hc0;
      11'd214  : in_data <= 8'h1c;
      11'd215  : in_data <= 8'hfd;
      11'd216  : in_data <= 8'ha3;
      11'd217  : in_data <= 8'h55;
      11'd218  : in_data <= 8'hf5;
      11'd219  : in_data <= 8'h77;
      11'd220  : in_data <= 8'h05;
      11'd221  : in_data <= 8'heb;
      11'd222  : in_data <= 8'hcb;
      11'd223  : in_data <= 8'he3;
      11'd224  : in_data <= 8'h9c;
      11'd225  : in_data <= 8'h4d;
      11'd226  : in_data <= 8'h13;
      11'd227  : in_data <= 8'hef;
      11'd228  : in_data <= 8'h6b;
      11'd229  : in_data <= 8'h2f;
      11'd230  : in_data <= 8'hba;
      11'd231  : in_data <= 8'h94;
      11'd232  : in_data <= 8'he0;
      11'd233  : in_data <= 8'h7a;
      11'd234  : in_data <= 8'h97;
      11'd235  : in_data <= 8'h35;
      11'd236  : in_data <= 8'h5d;
      11'd237  : in_data <= 8'h0e;
      11'd238  : in_data <= 8'h2a;
      11'd239  : in_data <= 8'h4c;
      11'd240  : in_data <= 8'hc9;
      11'd241  : in_data <= 8'hd7;
      11'd242  : in_data <= 8'h7e;
      11'd243  : in_data <= 8'h56;
      11'd244  : in_data <= 8'h85;
      11'd245  : in_data <= 8'h62;
      11'd246  : in_data <= 8'h23;
      11'd247  : in_data <= 8'hbe;
      11'd248  : in_data <= 8'h6c;
      11'd249  : in_data <= 8'hda;
      11'd250  : in_data <= 8'h04;
      11'd251  : in_data <= 8'hb0;
      11'd252  : in_data <= 8'hd9;
      11'd253  : in_data <= 8'h31;
      11'd254  : in_data <= 8'h04;
      11'd255  : in_data <= 8'h3f;
      11'd256  : in_data <= 8'hb0;
      11'd257  : in_data <= 8'h89;
      11'd258  : in_data <= 8'hc1;
      11'd259  : in_data <= 8'h6a;
      11'd260  : in_data <= 8'h1e;
      11'd261  : in_data <= 8'h69;
      11'd262  : in_data <= 8'hf0;
      11'd263  : in_data <= 8'hbe;
      11'd264  : in_data <= 8'hbc;
      11'd265  : in_data <= 8'h60;
      11'd266  : in_data <= 8'h1e;
      11'd267  : in_data <= 8'h7e;
      11'd268  : in_data <= 8'h42;
      11'd269  : in_data <= 8'hef;
      11'd270  : in_data <= 8'ha9;
      11'd271  : in_data <= 8'h45;
      11'd272  : in_data <= 8'hba;
      11'd273  : in_data <= 8'h0c;
      11'd274  : in_data <= 8'h5a;
      11'd275  : in_data <= 8'h20;
      11'd276  : in_data <= 8'he8;
      11'd277  : in_data <= 8'h46;
      11'd278  : in_data <= 8'ha2;
      11'd279  : in_data <= 8'h3a;
      11'd280  : in_data <= 8'h3d;
      11'd281  : in_data <= 8'h55;
      11'd282  : in_data <= 8'haa;
      11'd283  : in_data <= 8'hb1;
      11'd284  : in_data <= 8'hae;
      11'd285  : in_data <= 8'hb2;
      11'd286  : in_data <= 8'hcc;
      11'd287  : in_data <= 8'hdc;
      11'd288  : in_data <= 8'h85;
      11'd289  : in_data <= 8'h2e;
      11'd290  : in_data <= 8'he0;
      11'd291  : in_data <= 8'h16;
      11'd292  : in_data <= 8'h7b;
      11'd293  : in_data <= 8'h46;
      11'd294  : in_data <= 8'h93;
      11'd295  : in_data <= 8'h7d;
      11'd296  : in_data <= 8'h55;
      11'd297  : in_data <= 8'h9b;
      11'd298  : in_data <= 8'hcd;
      11'd299  : in_data <= 8'hc5;
      11'd300  : in_data <= 8'h27;
      11'd301  : in_data <= 8'hb2;
      11'd302  : in_data <= 8'h09;
      11'd303  : in_data <= 8'h50;
      11'd304  : in_data <= 8'h99;
      11'd305  : in_data <= 8'h1e;
      11'd306  : in_data <= 8'hef;
      11'd307  : in_data <= 8'h22;
      11'd308  : in_data <= 8'he0;
      11'd309  : in_data <= 8'ha9;
      11'd310  : in_data <= 8'hdc;
      11'd311  : in_data <= 8'h24;
      11'd312  : in_data <= 8'h18;
      11'd313  : in_data <= 8'hf4;
      11'd314  : in_data <= 8'hbc;
      11'd315  : in_data <= 8'h51;
      11'd316  : in_data <= 8'h8f;
      11'd317  : in_data <= 8'h4c;
      11'd318  : in_data <= 8'ha1;
      11'd319  : in_data <= 8'h1b;
      11'd320  : in_data <= 8'h5d;
      11'd321  : in_data <= 8'hba;
      11'd322  : in_data <= 8'h5a;
      11'd323  : in_data <= 8'h9b;
      11'd324  : in_data <= 8'hb2;
      11'd325  : in_data <= 8'hc9;
      11'd326  : in_data <= 8'h8f;
      11'd327  : in_data <= 8'hc5;
      11'd328  : in_data <= 8'hb1;
      11'd329  : in_data <= 8'h14;
      11'd330  : in_data <= 8'h4c;
      11'd331  : in_data <= 8'h36;
      11'd332  : in_data <= 8'h70;
      11'd333  : in_data <= 8'hdd;
      11'd334  : in_data <= 8'h60;
      11'd335  : in_data <= 8'h5c;
      11'd336  : in_data <= 8'h76;
      11'd337  : in_data <= 8'hcf;
      11'd338  : in_data <= 8'h51;
      11'd339  : in_data <= 8'h4f;
      11'd340  : in_data <= 8'h82;
      11'd341  : in_data <= 8'h0d;
      11'd342  : in_data <= 8'hcc;
      11'd343  : in_data <= 8'hae;
      11'd344  : in_data <= 8'h4b;
      11'd345  : in_data <= 8'h8b;
      11'd346  : in_data <= 8'h17;
      11'd347  : in_data <= 8'h8b;
      11'd348  : in_data <= 8'h27;
      11'd349  : in_data <= 8'hd1;
      11'd350  : in_data <= 8'heb;
      11'd351  : in_data <= 8'h04;
      11'd352  : in_data <= 8'h09;
      11'd353  : in_data <= 8'hbe;
      11'd354  : in_data <= 8'h0d;
      11'd355  : in_data <= 8'h1c;
      11'd356  : in_data <= 8'h14;
      11'd357  : in_data <= 8'h39;
      11'd358  : in_data <= 8'hc6;
      11'd359  : in_data <= 8'h69;
      11'd360  : in_data <= 8'hc7;
      11'd361  : in_data <= 8'hb5;
      11'd362  : in_data <= 8'h53;
      11'd363  : in_data <= 8'hec;
      11'd364  : in_data <= 8'h1d;
      11'd365  : in_data <= 8'hbf;
      11'd366  : in_data <= 8'h41;
      11'd367  : in_data <= 8'h58;
      11'd368  : in_data <= 8'hc8;
      11'd369  : in_data <= 8'h00;
      11'd370  : in_data <= 8'h69;
      11'd371  : in_data <= 8'h52;
      11'd372  : in_data <= 8'h09;
      11'd373  : in_data <= 8'h2f;
      11'd374  : in_data <= 8'hf0;
      11'd375  : in_data <= 8'h2f;
      11'd376  : in_data <= 8'hdd;
      11'd377  : in_data <= 8'ha5;
      11'd378  : in_data <= 8'h1c;
      11'd379  : in_data <= 8'ha0;
      11'd380  : in_data <= 8'h57;
      11'd381  : in_data <= 8'hae;
      11'd382  : in_data <= 8'h2f;
      11'd383  : in_data <= 8'h96;
      11'd384  : in_data <= 8'h82;
      11'd385  : in_data <= 8'ha4;
      11'd386  : in_data <= 8'h4b;
      11'd387  : in_data <= 8'h85;
      11'd388  : in_data <= 8'hd6;
      11'd389  : in_data <= 8'hab;
      11'd390  : in_data <= 8'hf4;
      11'd391  : in_data <= 8'h1f;
      11'd392  : in_data <= 8'h7b;
      11'd393  : in_data <= 8'hc5;
      11'd394  : in_data <= 8'h94;
      11'd395  : in_data <= 8'h1a;
      11'd396  : in_data <= 8'h73;
      11'd397  : in_data <= 8'h2d;
      11'd398  : in_data <= 8'h3a;
      11'd399  : in_data <= 8'h38;
      11'd400  : in_data <= 8'hea;
      11'd401  : in_data <= 8'hfc;
      11'd402  : in_data <= 8'hff;
      11'd403  : in_data <= 8'h81;
      11'd404  : in_data <= 8'h52;
      11'd405  : in_data <= 8'h06;
      11'd406  : in_data <= 8'h49;
      11'd407  : in_data <= 8'hd5;
      11'd408  : in_data <= 8'h97;
      11'd409  : in_data <= 8'hb4;
      11'd410  : in_data <= 8'h8b;
      11'd411  : in_data <= 8'ha2;
      11'd412  : in_data <= 8'h9e;
      11'd413  : in_data <= 8'h44;
      11'd414  : in_data <= 8'hcf;
      11'd415  : in_data <= 8'hb0;
      11'd416  : in_data <= 8'h8c;
      11'd417  : in_data <= 8'h4b;
      11'd418  : in_data <= 8'hd5;
      11'd419  : in_data <= 8'h82;
      11'd420  : in_data <= 8'h4d;
      11'd421  : in_data <= 8'h8a;
      11'd422  : in_data <= 8'hf4;
      11'd423  : in_data <= 8'h7a;
      11'd424  : in_data <= 8'h85;
      11'd425  : in_data <= 8'hee;
      11'd426  : in_data <= 8'hfe;
      11'd427  : in_data <= 8'hd0;
      11'd428  : in_data <= 8'h25;
      11'd429  : in_data <= 8'h9c;
      11'd430  : in_data <= 8'h7a;
      11'd431  : in_data <= 8'h4a;
      11'd432  : in_data <= 8'h57;
      11'd433  : in_data <= 8'hf6;
      11'd434  : in_data <= 8'h8b;
      11'd435  : in_data <= 8'hf7;
      11'd436  : in_data <= 8'h09;
      11'd437  : in_data <= 8'ha3;
      11'd438  : in_data <= 8'h27;
      11'd439  : in_data <= 8'h74;
      11'd440  : in_data <= 8'h31;
      11'd441  : in_data <= 8'had;
      11'd442  : in_data <= 8'h87;
      11'd443  : in_data <= 8'hda;
      11'd444  : in_data <= 8'h13;
      11'd445  : in_data <= 8'hf2;
      11'd446  : in_data <= 8'h81;
      11'd447  : in_data <= 8'h1e;
      11'd448  : in_data <= 8'h78;
      11'd449  : in_data <= 8'h83;
      11'd450  : in_data <= 8'h34;
      11'd451  : in_data <= 8'he1;
      11'd452  : in_data <= 8'h83;
      11'd453  : in_data <= 8'h46;
      11'd454  : in_data <= 8'hde;
      11'd455  : in_data <= 8'h6f;
      11'd456  : in_data <= 8'h82;
      11'd457  : in_data <= 8'h22;
      11'd458  : in_data <= 8'h74;
      11'd459  : in_data <= 8'h6a;
      11'd460  : in_data <= 8'h39;
      11'd461  : in_data <= 8'hc6;
      11'd462  : in_data <= 8'h00;
      11'd463  : in_data <= 8'hfd;
      11'd464  : in_data <= 8'hdc;
      11'd465  : in_data <= 8'hfd;
      11'd466  : in_data <= 8'he5;
      11'd467  : in_data <= 8'h9d;
      11'd468  : in_data <= 8'hc9;
      11'd469  : in_data <= 8'h86;
      11'd470  : in_data <= 8'h1c;
      11'd471  : in_data <= 8'h8d;
      11'd472  : in_data <= 8'h0e;
      11'd473  : in_data <= 8'h09;
      11'd474  : in_data <= 8'h5a;
      11'd475  : in_data <= 8'he2;
      11'd476  : in_data <= 8'h6d;
      11'd477  : in_data <= 8'h26;
      11'd478  : in_data <= 8'hd3;
      11'd479  : in_data <= 8'ha8;
      11'd480  : in_data <= 8'h28;
      11'd481  : in_data <= 8'h11;
      11'd482  : in_data <= 8'h1a;
      11'd483  : in_data <= 8'h36;
      11'd484  : in_data <= 8'hf2;
      11'd485  : in_data <= 8'h93;
      11'd486  : in_data <= 8'he0;
      11'd487  : in_data <= 8'h73;
      11'd488  : in_data <= 8'h37;
      11'd489  : in_data <= 8'h57;
      11'd490  : in_data <= 8'hdd;
      11'd491  : in_data <= 8'h35;
      11'd492  : in_data <= 8'hfa;
      11'd493  : in_data <= 8'h5d;
      11'd494  : in_data <= 8'hbd;
      11'd495  : in_data <= 8'h6a;
      11'd496  : in_data <= 8'h7d;
      11'd497  : in_data <= 8'h0a;
      11'd498  : in_data <= 8'h81;
      11'd499  : in_data <= 8'hda;
      11'd500  : in_data <= 8'h9e;
      11'd501  : in_data <= 8'h8c;
      11'd502  : in_data <= 8'h26;
      11'd503  : in_data <= 8'h53;
      11'd504  : in_data <= 8'h5c;
      11'd505  : in_data <= 8'hf3;
      11'd506  : in_data <= 8'hd7;
      11'd507  : in_data <= 8'h7a;
      11'd508  : in_data <= 8'h26;
      11'd509  : in_data <= 8'h26;
      11'd510  : in_data <= 8'hfb;
      11'd511  : in_data <= 8'hf2;
      11'd512  : in_data <= 8'ha4;
      11'd513  : in_data <= 8'hf3;
      11'd514  : in_data <= 8'h19;
      11'd515  : in_data <= 8'h70;
      11'd516  : in_data <= 8'hf4;
      11'd517  : in_data <= 8'h8d;
      11'd518  : in_data <= 8'h05;
      11'd519  : in_data <= 8'hfe;
      11'd520  : in_data <= 8'h57;
      11'd521  : in_data <= 8'h58;
      11'd522  : in_data <= 8'hfd;
      11'd523  : in_data <= 8'h0e;
      11'd524  : in_data <= 8'hb8;
      11'd525  : in_data <= 8'hf7;
      11'd526  : in_data <= 8'hbb;
      11'd527  : in_data <= 8'haa;
      11'd528  : in_data <= 8'h76;
      11'd529  : in_data <= 8'h7b;
      11'd530  : in_data <= 8'hf8;
      11'd531  : in_data <= 8'h61;
      11'd532  : in_data <= 8'hd6;
      11'd533  : in_data <= 8'h85;
      11'd534  : in_data <= 8'h69;
      11'd535  : in_data <= 8'hea;
      11'd536  : in_data <= 8'haf;
      11'd537  : in_data <= 8'h23;
      11'd538  : in_data <= 8'h10;
      11'd539  : in_data <= 8'h48;
      11'd540  : in_data <= 8'h02;
      11'd541  : in_data <= 8'h11;
      11'd542  : in_data <= 8'h12;
      11'd543  : in_data <= 8'hc8;
      11'd544  : in_data <= 8'h54;
      11'd545  : in_data <= 8'h5e;
      11'd546  : in_data <= 8'h15;
      11'd547  : in_data <= 8'h88;
      11'd548  : in_data <= 8'h32;
      11'd549  : in_data <= 8'he0;
      11'd550  : in_data <= 8'h02;
      11'd551  : in_data <= 8'h5e;
      11'd552  : in_data <= 8'h57;
      11'd553  : in_data <= 8'hb7;
      11'd554  : in_data <= 8'hd6;
      11'd555  : in_data <= 8'h47;
      11'd556  : in_data <= 8'h6f;
      11'd557  : in_data <= 8'h01;
      11'd558  : in_data <= 8'heb;
      11'd559  : in_data <= 8'h1b;
      11'd560  : in_data <= 8'h91;
      11'd561  : in_data <= 8'hb1;
      11'd562  : in_data <= 8'h1c;
      11'd563  : in_data <= 8'ha1;
      11'd564  : in_data <= 8'hd7;
      11'd565  : in_data <= 8'h2e;
      11'd566  : in_data <= 8'h57;
      11'd567  : in_data <= 8'hae;
      11'd568  : in_data <= 8'h46;
      11'd569  : in_data <= 8'h82;
      11'd570  : in_data <= 8'h86;
      11'd571  : in_data <= 8'h12;
      11'd572  : in_data <= 8'h52;
      11'd573  : in_data <= 8'he0;
      11'd574  : in_data <= 8'hfd;
      11'd575  : in_data <= 8'ha1;
      11'd576  : in_data <= 8'hb6;
      11'd577  : in_data <= 8'hc0;
      11'd578  : in_data <= 8'hfb;
      11'd579  : in_data <= 8'h59;
      11'd580  : in_data <= 8'hf9;
      11'd581  : in_data <= 8'h10;
      11'd582  : in_data <= 8'h15;
      11'd583  : in_data <= 8'h76;
      11'd584  : in_data <= 8'h3a;
      11'd585  : in_data <= 8'h38;
      11'd586  : in_data <= 8'h7b;
      11'd587  : in_data <= 8'hbd;
      11'd588  : in_data <= 8'he6;
      11'd589  : in_data <= 8'h11;
      11'd590  : in_data <= 8'h9a;
      11'd591  : in_data <= 8'h59;
      11'd592  : in_data <= 8'hd0;
      11'd593  : in_data <= 8'h87;
      11'd594  : in_data <= 8'h92;
      11'd595  : in_data <= 8'hef;
      11'd596  : in_data <= 8'hcd;
      11'd597  : in_data <= 8'hf5;
      11'd598  : in_data <= 8'h2e;
      11'd599  : in_data <= 8'had;
      11'd600  : in_data <= 8'h78;
      11'd601  : in_data <= 8'h01;
      11'd602  : in_data <= 8'h8b;
      11'd603  : in_data <= 8'h46;
      11'd604  : in_data <= 8'h34;
      11'd605  : in_data <= 8'hbb;
      11'd606  : in_data <= 8'h65;
      11'd607  : in_data <= 8'hbc;
      11'd608  : in_data <= 8'h9d;
      11'd609  : in_data <= 8'h97;
      11'd610  : in_data <= 8'hf3;
      11'd611  : in_data <= 8'h6c;
      11'd612  : in_data <= 8'hc8;
      11'd613  : in_data <= 8'h89;
      11'd614  : in_data <= 8'he6;
      11'd615  : in_data <= 8'hb9;
      11'd616  : in_data <= 8'h8f;
      11'd617  : in_data <= 8'h15;
      11'd618  : in_data <= 8'h2f;
      11'd619  : in_data <= 8'h61;
      11'd620  : in_data <= 8'hf2;
      11'd621  : in_data <= 8'h42;
      11'd622  : in_data <= 8'h35;
      11'd623  : in_data <= 8'h36;
      11'd624  : in_data <= 8'h55;
      11'd625  : in_data <= 8'ha4;
      11'd626  : in_data <= 8'hb2;
      11'd627  : in_data <= 8'h30;
      11'd628  : in_data <= 8'h1b;
      11'd629  : in_data <= 8'hd4;
      11'd630  : in_data <= 8'h46;
      11'd631  : in_data <= 8'h5a;
      11'd632  : in_data <= 8'h68;
      11'd633  : in_data <= 8'hff;
      11'd634  : in_data <= 8'h61;
      11'd635  : in_data <= 8'h67;
      11'd636  : in_data <= 8'he0;
      11'd637  : in_data <= 8'ha7;
      11'd638  : in_data <= 8'ha8;
      11'd639  : in_data <= 8'h4d;
      11'd640  : in_data <= 8'h7b;
      11'd641  : in_data <= 8'hec;
      11'd642  : in_data <= 8'ha4;
      11'd643  : in_data <= 8'ha3;
      11'd644  : in_data <= 8'h1a;
      11'd645  : in_data <= 8'h43;
      11'd646  : in_data <= 8'h93;
      11'd647  : in_data <= 8'h18;
      11'd648  : in_data <= 8'h2b;
      11'd649  : in_data <= 8'hd7;
      11'd650  : in_data <= 8'h74;
      11'd651  : in_data <= 8'h0e;
      11'd652  : in_data <= 8'h6b;
      11'd653  : in_data <= 8'hf9;
      11'd654  : in_data <= 8'h3d;
      11'd655  : in_data <= 8'hf0;
      11'd656  : in_data <= 8'he9;
      11'd657  : in_data <= 8'hbf;
      11'd658  : in_data <= 8'h7a;
      11'd659  : in_data <= 8'h72;
      11'd660  : in_data <= 8'h5e;
      11'd661  : in_data <= 8'h1d;
      11'd662  : in_data <= 8'heb;
      11'd663  : in_data <= 8'he7;
      11'd664  : in_data <= 8'h92;
      11'd665  : in_data <= 8'h4d;
      11'd666  : in_data <= 8'h2e;
      11'd667  : in_data <= 8'h93;
      11'd668  : in_data <= 8'hfc;
      11'd669  : in_data <= 8'h1c;
      11'd670  : in_data <= 8'ha9;
      11'd671  : in_data <= 8'h3e;
      11'd672  : in_data <= 8'h2a;
      11'd673  : in_data <= 8'h1f;
      11'd674  : in_data <= 8'hb7;
      11'd675  : in_data <= 8'hf6;
      11'd676  : in_data <= 8'h78;
      11'd677  : in_data <= 8'h4e;
      11'd678  : in_data <= 8'h70;
      11'd679  : in_data <= 8'hcf;
      11'd680  : in_data <= 8'h22;
      11'd681  : in_data <= 8'ha8;
      11'd682  : in_data <= 8'h18;
      11'd683  : in_data <= 8'hb1;
      11'd684  : in_data <= 8'h74;
      11'd685  : in_data <= 8'h78;
      11'd686  : in_data <= 8'h40;
      11'd687  : in_data <= 8'hfe;
      11'd688  : in_data <= 8'ha8;
      11'd689  : in_data <= 8'hfd;
      11'd690  : in_data <= 8'h5d;
      11'd691  : in_data <= 8'h59;
      11'd692  : in_data <= 8'h82;
      11'd693  : in_data <= 8'hff;
      11'd694  : in_data <= 8'h1e;
      11'd695  : in_data <= 8'h63;
      11'd696  : in_data <= 8'hcc;
      11'd697  : in_data <= 8'h46;
      11'd698  : in_data <= 8'h63;
      11'd699  : in_data <= 8'h50;
      11'd700  : in_data <= 8'h21;
      11'd701  : in_data <= 8'h57;
      11'd702  : in_data <= 8'h18;
      11'd703  : in_data <= 8'h46;
      11'd704  : in_data <= 8'h5a;
      11'd705  : in_data <= 8'h50;
      11'd706  : in_data <= 8'h11;
      11'd707  : in_data <= 8'h9c;
      11'd708  : in_data <= 8'h95;
      11'd709  : in_data <= 8'hb1;
      11'd710  : in_data <= 8'h11;
      11'd711  : in_data <= 8'hc6;
      11'd712  : in_data <= 8'hc7;
      11'd713  : in_data <= 8'h6d;
      11'd714  : in_data <= 8'h97;
      11'd715  : in_data <= 8'h5b;
      11'd716  : in_data <= 8'h71;
      11'd717  : in_data <= 8'h2d;
      11'd718  : in_data <= 8'hf9;
      11'd719  : in_data <= 8'h27;
      11'd720  : in_data <= 8'h46;
      11'd721  : in_data <= 8'h56;
      11'd722  : in_data <= 8'hf6;
      11'd723  : in_data <= 8'h0f;
      11'd724  : in_data <= 8'h2e;
      11'd725  : in_data <= 8'h16;
      11'd726  : in_data <= 8'h86;
      11'd727  : in_data <= 8'hbb;
      11'd728  : in_data <= 8'h8d;
      11'd729  : in_data <= 8'h01;
      11'd730  : in_data <= 8'h7e;
      11'd731  : in_data <= 8'h10;
      11'd732  : in_data <= 8'h2a;
      11'd733  : in_data <= 8'h94;
      11'd734  : in_data <= 8'h7e;
      11'd735  : in_data <= 8'hf4;
      11'd736  : in_data <= 8'hef;
      11'd737  : in_data <= 8'h9b;
      11'd738  : in_data <= 8'h6f;
      11'd739  : in_data <= 8'hd7;
      11'd740  : in_data <= 8'hf3;
      11'd741  : in_data <= 8'hed;
      11'd742  : in_data <= 8'ha0;
      11'd743  : in_data <= 8'he2;
      11'd744  : in_data <= 8'hbb;
      11'd745  : in_data <= 8'hd6;
      11'd746  : in_data <= 8'h42;
      11'd747  : in_data <= 8'h4b;
      11'd748  : in_data <= 8'h24;
      11'd749  : in_data <= 8'hf8;
      11'd750  : in_data <= 8'h02;
      11'd751  : in_data <= 8'h7c;
      11'd752  : in_data <= 8'h7a;
      11'd753  : in_data <= 8'h60;
      11'd754  : in_data <= 8'ha4;
      11'd755  : in_data <= 8'h3a;
      11'd756  : in_data <= 8'hb5;
      11'd757  : in_data <= 8'h1a;
      11'd758  : in_data <= 8'h7c;
      11'd759  : in_data <= 8'h94;
      11'd760  : in_data <= 8'hdd;
      11'd761  : in_data <= 8'hbb;
      11'd762  : in_data <= 8'h96;
      11'd763  : in_data <= 8'h81;
      11'd764  : in_data <= 8'he0;
      11'd765  : in_data <= 8'h33;
      11'd766  : in_data <= 8'hf4;
      11'd767  : in_data <= 8'h9b;
      11'd768  : in_data <= 8'h54;
      11'd769  : in_data <= 8'h13;
      11'd770  : in_data <= 8'h02;
      11'd771  : in_data <= 8'ha3;
      11'd772  : in_data <= 8'h66;
      11'd773  : in_data <= 8'h79;
      11'd774  : in_data <= 8'h76;
      11'd775  : in_data <= 8'h4e;
      11'd776  : in_data <= 8'ha3;
      11'd777  : in_data <= 8'h7d;
      11'd778  : in_data <= 8'hc4;
      11'd779  : in_data <= 8'h4f;
      11'd780  : in_data <= 8'h23;
      11'd781  : in_data <= 8'h93;
      11'd782  : in_data <= 8'h22;
      11'd783  : in_data <= 8'h3c;
      11'd784  : in_data <= 8'h78;
      11'd785  : in_data <= 8'h72;
      11'd786  : in_data <= 8'h8b;
      11'd787  : in_data <= 8'hb8;
      11'd788  : in_data <= 8'hcc;
      11'd789  : in_data <= 8'ha6;
      11'd790  : in_data <= 8'h9f;
      11'd791  : in_data <= 8'had;
      11'd792  : in_data <= 8'hfa;
      11'd793  : in_data <= 8'ha6;
      11'd794  : in_data <= 8'hdf;
      11'd795  : in_data <= 8'hc6;
      11'd796  : in_data <= 8'hd1;
      11'd797  : in_data <= 8'h7f;
      11'd798  : in_data <= 8'h96;
      11'd799  : in_data <= 8'h8b;
      11'd800  : in_data <= 8'hfd;
      11'd801  : in_data <= 8'h1d;
      11'd802  : in_data <= 8'h45;
      11'd803  : in_data <= 8'h24;
      11'd804  : in_data <= 8'h52;
      11'd805  : in_data <= 8'hf0;
      11'd806  : in_data <= 8'hca;
      11'd807  : in_data <= 8'h4d;
      11'd808  : in_data <= 8'ha9;
      11'd809  : in_data <= 8'hfd;
      11'd810  : in_data <= 8'h3e;
      11'd811  : in_data <= 8'h67;
      11'd812  : in_data <= 8'hbe;
      11'd813  : in_data <= 8'hd7;
      11'd814  : in_data <= 8'h82;
      11'd815  : in_data <= 8'hdc;
      11'd816  : in_data <= 8'hd6;
      11'd817  : in_data <= 8'h40;
      11'd818  : in_data <= 8'h02;
      11'd819  : in_data <= 8'h35;
      11'd820  : in_data <= 8'h44;
      11'd821  : in_data <= 8'h2f;
      11'd822  : in_data <= 8'haa;
      11'd823  : in_data <= 8'h8d;
      11'd824  : in_data <= 8'h42;
      11'd825  : in_data <= 8'h93;
      11'd826  : in_data <= 8'h76;
      11'd827  : in_data <= 8'h7b;
      11'd828  : in_data <= 8'he7;
      11'd829  : in_data <= 8'hc9;
      11'd830  : in_data <= 8'h1f;
      11'd831  : in_data <= 8'hdc;
      11'd832  : in_data <= 8'h74;
      11'd833  : in_data <= 8'h3d;
      11'd834  : in_data <= 8'hba;
      11'd835  : in_data <= 8'h9b;
      11'd836  : in_data <= 8'hfe;
      11'd837  : in_data <= 8'h59;
      11'd838  : in_data <= 8'h10;
      11'd839  : in_data <= 8'h67;
      11'd840  : in_data <= 8'h47;
      11'd841  : in_data <= 8'h49;
      11'd842  : in_data <= 8'ha1;
      11'd843  : in_data <= 8'hb1;
      11'd844  : in_data <= 8'hfa;
      11'd845  : in_data <= 8'h5c;
      11'd846  : in_data <= 8'hb3;
      11'd847  : in_data <= 8'h38;
      11'd848  : in_data <= 8'h10;
      11'd849  : in_data <= 8'h6f;
      11'd850  : in_data <= 8'hb3;
      11'd851  : in_data <= 8'h82;
      11'd852  : in_data <= 8'h8d;
      11'd853  : in_data <= 8'h0c;
      11'd854  : in_data <= 8'ha7;
      11'd855  : in_data <= 8'h32;
      11'd856  : in_data <= 8'h03;
      11'd857  : in_data <= 8'h77;
      11'd858  : in_data <= 8'h00;
      11'd859  : in_data <= 8'h35;
      11'd860  : in_data <= 8'h51;
      11'd861  : in_data <= 8'h8d;
      11'd862  : in_data <= 8'hfa;
      11'd863  : in_data <= 8'h4b;
      11'd864  : in_data <= 8'h92;
      11'd865  : in_data <= 8'h0f;
      11'd866  : in_data <= 8'hc2;
      11'd867  : in_data <= 8'hfa;
      11'd868  : in_data <= 8'heb;
      11'd869  : in_data <= 8'h2a;
      11'd870  : in_data <= 8'h1c;
      11'd871  : in_data <= 8'h99;
      11'd872  : in_data <= 8'hf4;
      11'd873  : in_data <= 8'hb6;
      11'd874  : in_data <= 8'he0;
      11'd875  : in_data <= 8'h39;
      11'd876  : in_data <= 8'h3f;
      11'd877  : in_data <= 8'h9b;
      11'd878  : in_data <= 8'hbb;
      11'd879  : in_data <= 8'h00;
      11'd880  : in_data <= 8'h9c;
      11'd881  : in_data <= 8'h64;
      11'd882  : in_data <= 8'ha2;
      11'd883  : in_data <= 8'h1c;
      11'd884  : in_data <= 8'h43;
      11'd885  : in_data <= 8'h17;
      11'd886  : in_data <= 8'hf6;
      11'd887  : in_data <= 8'h2f;
      11'd888  : in_data <= 8'h7f;
      11'd889  : in_data <= 8'h0b;
      11'd890  : in_data <= 8'h00;
      11'd891  : in_data <= 8'h20;
      11'd892  : in_data <= 8'h18;
      11'd893  : in_data <= 8'hb0;
      11'd894  : in_data <= 8'hfd;
      11'd895  : in_data <= 8'he4;
      11'd896  : in_data <= 8'h67;
      11'd897  : in_data <= 8'hc1;
      11'd898  : in_data <= 8'h4c;
      11'd899  : in_data <= 8'hf8;
      11'd900  : in_data <= 8'h68;
      11'd901  : in_data <= 8'h48;
      11'd902  : in_data <= 8'h30;
      11'd903  : in_data <= 8'h4c;
      11'd904  : in_data <= 8'hc6;
      11'd905  : in_data <= 8'h32;
      11'd906  : in_data <= 8'he0;
      11'd907  : in_data <= 8'h35;
      11'd908  : in_data <= 8'h62;
      11'd909  : in_data <= 8'ha7;
      11'd910  : in_data <= 8'h16;
      11'd911  : in_data <= 8'h94;
      11'd912  : in_data <= 8'h7a;
      11'd913  : in_data <= 8'h32;
      11'd914  : in_data <= 8'hb4;
      11'd915  : in_data <= 8'h23;
      11'd916  : in_data <= 8'h07;
      11'd917  : in_data <= 8'h99;
      11'd918  : in_data <= 8'h63;
      11'd919  : in_data <= 8'hfa;
      11'd920  : in_data <= 8'hfa;
      11'd921  : in_data <= 8'hd2;
      11'd922  : in_data <= 8'h96;
      11'd923  : in_data <= 8'he7;
      11'd924  : in_data <= 8'h81;
      11'd925  : in_data <= 8'h03;
      11'd926  : in_data <= 8'h08;
      11'd927  : in_data <= 8'h83;
      11'd928  : in_data <= 8'hd4;
      11'd929  : in_data <= 8'hc8;
      11'd930  : in_data <= 8'h29;
      11'd931  : in_data <= 8'h7b;
      11'd932  : in_data <= 8'h9c;
      11'd933  : in_data <= 8'h4d;
      11'd934  : in_data <= 8'h41;
      11'd935  : in_data <= 8'hfc;
      11'd936  : in_data <= 8'hcf;
      11'd937  : in_data <= 8'h86;
      11'd938  : in_data <= 8'hd9;
      11'd939  : in_data <= 8'h4b;
      11'd940  : in_data <= 8'hc4;
      11'd941  : in_data <= 8'h8a;
      11'd942  : in_data <= 8'hde;
      11'd943  : in_data <= 8'hfb;
      11'd944  : in_data <= 8'h11;
      11'd945  : in_data <= 8'ha3;
      11'd946  : in_data <= 8'hb9;
      11'd947  : in_data <= 8'h3a;
      11'd948  : in_data <= 8'h68;
      11'd949  : in_data <= 8'h76;
      11'd950  : in_data <= 8'h16;
      11'd951  : in_data <= 8'h14;
      11'd952  : in_data <= 8'h9f;
      11'd953  : in_data <= 8'hca;
      11'd954  : in_data <= 8'h1c;
      11'd955  : in_data <= 8'h44;
      11'd956  : in_data <= 8'ha7;
      11'd957  : in_data <= 8'hc6;
      11'd958  : in_data <= 8'h00;
      11'd959  : in_data <= 8'h16;
      11'd960  : in_data <= 8'h02;
      11'd961  : in_data <= 8'h59;
      11'd962  : in_data <= 8'hb2;
      11'd963  : in_data <= 8'h71;
      11'd964  : in_data <= 8'hfb;
      11'd965  : in_data <= 8'h41;
      11'd966  : in_data <= 8'h1c;
      11'd967  : in_data <= 8'hc9;
      11'd968  : in_data <= 8'hc5;
      11'd969  : in_data <= 8'h39;
      11'd970  : in_data <= 8'hf2;
      11'd971  : in_data <= 8'h54;
      11'd972  : in_data <= 8'haa;
      11'd973  : in_data <= 8'hc7;
      11'd974  : in_data <= 8'h1c;
      11'd975  : in_data <= 8'hd1;
      11'd976  : in_data <= 8'h93;
      11'd977  : in_data <= 8'ha6;
      11'd978  : in_data <= 8'h96;
      11'd979  : in_data <= 8'h23;
      11'd980  : in_data <= 8'h9f;
      11'd981  : in_data <= 8'h3c;
      11'd982  : in_data <= 8'h09;
      11'd983  : in_data <= 8'h99;
      11'd984  : in_data <= 8'h28;
      11'd985  : in_data <= 8'ha6;
      11'd986  : in_data <= 8'hbf;
      11'd987  : in_data <= 8'hca;
      11'd988  : in_data <= 8'hd5;
      11'd989  : in_data <= 8'h8b;
      11'd990  : in_data <= 8'h29;
      11'd991  : in_data <= 8'hd9;
      11'd992  : in_data <= 8'he9;
      11'd993  : in_data <= 8'hfe;
      11'd994  : in_data <= 8'h6a;
      11'd995  : in_data <= 8'h57;
      11'd996  : in_data <= 8'h36;
      11'd997  : in_data <= 8'h88;
      11'd998  : in_data <= 8'hac;
      11'd999  : in_data <= 8'had;
      11'd1000 : in_data <= 8'h23;
      11'd1001 : in_data <= 8'hbd;
      11'd1002 : in_data <= 8'h58;
      11'd1003 : in_data <= 8'h9a;
      11'd1004 : in_data <= 8'h19;
      11'd1005 : in_data <= 8'h51;
      11'd1006 : in_data <= 8'h1b;
      11'd1007 : in_data <= 8'h35;
      11'd1008 : in_data <= 8'h0b;
      11'd1009 : in_data <= 8'h70;
      11'd1010 : in_data <= 8'h26;
      11'd1011 : in_data <= 8'h78;
      11'd1012 : in_data <= 8'h1a;
      11'd1013 : in_data <= 8'h16;
      11'd1014 : in_data <= 8'h2b;
      11'd1015 : in_data <= 8'hac;
      11'd1016 : in_data <= 8'h46;
      11'd1017 : in_data <= 8'hb9;
      11'd1018 : in_data <= 8'h31;
      11'd1019 : in_data <= 8'hc6;
      11'd1020 : in_data <= 8'h85;
      11'd1021 : in_data <= 8'h61;
      11'd1022 : in_data <= 8'h86;
      11'd1023 : in_data <= 8'h4a;
      11'd1024 : in_data <= 8'h7b;
      11'd1025 : in_data <= 8'h9f;
      11'd1026 : in_data <= 8'hc1;
      11'd1027 : in_data <= 8'hff;
      11'd1028 : in_data <= 8'h32;
      11'd1029 : in_data <= 8'h4f;
      11'd1030 : in_data <= 8'h2d;
      11'd1031 : in_data <= 8'ha6;
      11'd1032 : in_data <= 8'h97;
      11'd1033 : in_data <= 8'hae;
      11'd1034 : in_data <= 8'h86;
      11'd1035 : in_data <= 8'ha0;
      11'd1036 : in_data <= 8'h75;
      11'd1037 : in_data <= 8'h5e;
      11'd1038 : in_data <= 8'h82;
      11'd1039 : in_data <= 8'h8e;
      11'd1040 : in_data <= 8'hb2;
      11'd1041 : in_data <= 8'h7e;
      11'd1042 : in_data <= 8'h3e;
      11'd1043 : in_data <= 8'h67;
      11'd1044 : in_data <= 8'h68;
      11'd1045 : in_data <= 8'h31;
      11'd1046 : in_data <= 8'h29;
      11'd1047 : in_data <= 8'h19;
      11'd1048 : in_data <= 8'h40;
      11'd1049 : in_data <= 8'h9f;
      11'd1050 : in_data <= 8'hfb;
      11'd1051 : in_data <= 8'h0b;
      11'd1052 : in_data <= 8'h19;
      11'd1053 : in_data <= 8'h25;
      11'd1054 : in_data <= 8'h8d;
      11'd1055 : in_data <= 8'h5b;
      11'd1056 : in_data <= 8'h72;
      11'd1057 : in_data <= 8'h9f;
      11'd1058 : in_data <= 8'h97;
      11'd1059 : in_data <= 8'hdf;
      11'd1060 : in_data <= 8'h43;
      11'd1061 : in_data <= 8'h39;
      11'd1062 : in_data <= 8'h99;
      11'd1063 : in_data <= 8'ha9;
      11'd1064 : in_data <= 8'hf9;
      11'd1065 : in_data <= 8'h55;
      11'd1066 : in_data <= 8'h38;
      11'd1067 : in_data <= 8'h16;
      11'd1068 : in_data <= 8'hd1;
      11'd1069 : in_data <= 8'h28;
      11'd1070 : in_data <= 8'h9a;
      11'd1071 : in_data <= 8'h62;
      11'd1072 : in_data <= 8'h07;
      11'd1073 : in_data <= 8'hc3;
      11'd1074 : in_data <= 8'h15;
      11'd1075 : in_data <= 8'hd8;
      11'd1076 : in_data <= 8'h1d;
      11'd1077 : in_data <= 8'hda;
      11'd1078 : in_data <= 8'h8e;
      11'd1079 : in_data <= 8'h57;
      11'd1080 : in_data <= 8'h13;
      11'd1081 : in_data <= 8'h96;
      11'd1082 : in_data <= 8'h6a;
      11'd1083 : in_data <= 8'hed;
      11'd1084 : in_data <= 8'h45;
      11'd1085 : in_data <= 8'hf9;
      11'd1086 : in_data <= 8'hec;
      11'd1087 : in_data <= 8'h7a;
      11'd1088 : in_data <= 8'h1b;
      11'd1089 : in_data <= 8'h24;
      11'd1090 : in_data <= 8'h59;
      11'd1091 : in_data <= 8'h2a;
      11'd1092 : in_data <= 8'h39;
      11'd1093 : in_data <= 8'h4c;
      11'd1094 : in_data <= 8'hdb;
      11'd1095 : in_data <= 8'ha3;
      11'd1096 : in_data <= 8'h7a;
      11'd1097 : in_data <= 8'h68;
      11'd1098 : in_data <= 8'he1;
      11'd1099 : in_data <= 8'had;
      11'd1100 : in_data <= 8'h9f;
      11'd1101 : in_data <= 8'h8a;
      11'd1102 : in_data <= 8'hdd;
      11'd1103 : in_data <= 8'h15;
      11'd1104 : in_data <= 8'h8e;
      11'd1105 : in_data <= 8'hf6;
      11'd1106 : in_data <= 8'h2c;
      11'd1107 : in_data <= 8'hf1;
      11'd1108 : in_data <= 8'h35;
      11'd1109 : in_data <= 8'h0c;
      11'd1110 : in_data <= 8'h37;
      11'd1111 : in_data <= 8'h03;
      11'd1112 : in_data <= 8'h25;
      11'd1113 : in_data <= 8'he0;
      11'd1114 : in_data <= 8'hf9;
      11'd1115 : in_data <= 8'hbe;
      11'd1116 : in_data <= 8'h61;
      11'd1117 : in_data <= 8'h5e;
      11'd1118 : in_data <= 8'h2c;
      11'd1119 : in_data <= 8'hf5;
      11'd1120 : in_data <= 8'hf5;
      11'd1121 : in_data <= 8'he1;
      11'd1122 : in_data <= 8'h9b;
      11'd1123 : in_data <= 8'h2c;
      11'd1124 : in_data <= 8'hc4;
      11'd1125 : in_data <= 8'he1;
      11'd1126 : in_data <= 8'h38;
      11'd1127 : in_data <= 8'h1e;
      11'd1128 : in_data <= 8'h25;
      11'd1129 : in_data <= 8'hd8;
      11'd1130 : in_data <= 8'hd1;
      11'd1131 : in_data <= 8'ha9;
      11'd1132 : in_data <= 8'h71;
      11'd1133 : in_data <= 8'h6c;
      11'd1134 : in_data <= 8'h8f;
      11'd1135 : in_data <= 8'h80;
      11'd1136 : in_data <= 8'hed;
      11'd1137 : in_data <= 8'hb7;
      11'd1138 : in_data <= 8'hf7;
      11'd1139 : in_data <= 8'h45;
      11'd1140 : in_data <= 8'h10;
      11'd1141 : in_data <= 8'h7c;
      11'd1142 : in_data <= 8'h68;
      11'd1143 : in_data <= 8'h81;
      11'd1144 : in_data <= 8'ha1;
      11'd1145 : in_data <= 8'hc2;
      11'd1146 : in_data <= 8'h05;
      11'd1147 : in_data <= 8'hde;
      11'd1148 : in_data <= 8'hab;
      11'd1149 : in_data <= 8'h59;
      11'd1150 : in_data <= 8'h37;
      11'd1151 : in_data <= 8'hba;
      11'd1152 : in_data <= 8'h6b;
      11'd1153 : in_data <= 8'hb7;
      11'd1154 : in_data <= 8'h87;
      11'd1155 : in_data <= 8'hc1;
      11'd1156 : in_data <= 8'h08;
      11'd1157 : in_data <= 8'h5c;
      11'd1158 : in_data <= 8'h6e;
      11'd1159 : in_data <= 8'h74;
      11'd1160 : in_data <= 8'hc8;
      11'd1161 : in_data <= 8'h2e;
      11'd1162 : in_data <= 8'h22;
      11'd1163 : in_data <= 8'h31;
      11'd1164 : in_data <= 8'h2f;
      11'd1165 : in_data <= 8'h80;
      11'd1166 : in_data <= 8'h9e;
      11'd1167 : in_data <= 8'h7a;
      11'd1168 : in_data <= 8'hb2;
      11'd1169 : in_data <= 8'h86;
      11'd1170 : in_data <= 8'he2;
      11'd1171 : in_data <= 8'h93;
      11'd1172 : in_data <= 8'ha4;
      11'd1173 : in_data <= 8'h07;
      11'd1174 : in_data <= 8'hf6;
      11'd1175 : in_data <= 8'hb2;
      11'd1176 : in_data <= 8'hf2;
      11'd1177 : in_data <= 8'h92;
      11'd1178 : in_data <= 8'hbe;
      11'd1179 : in_data <= 8'h0e;
      11'd1180 : in_data <= 8'hf0;
      11'd1181 : in_data <= 8'h4a;
      11'd1182 : in_data <= 8'hf6;
      11'd1183 : in_data <= 8'he6;
      11'd1184 : in_data <= 8'h9f;
      11'd1185 : in_data <= 8'h8b;
      11'd1186 : in_data <= 8'h37;
      11'd1187 : in_data <= 8'h50;
      11'd1188 : in_data <= 8'h0d;
      11'd1189 : in_data <= 8'ha3;
      11'd1190 : in_data <= 8'hd4;
      11'd1191 : in_data <= 8'h19;
      11'd1192 : in_data <= 8'heb;
      11'd1193 : in_data <= 8'hc8;
      11'd1194 : in_data <= 8'h72;
      11'd1195 : in_data <= 8'hc7;
      11'd1196 : in_data <= 8'he3;
      11'd1197 : in_data <= 8'h8f;
      11'd1198 : in_data <= 8'h59;
      11'd1199 : in_data <= 8'h7d;
      11'd1200 : in_data <= 8'h6f;
      11'd1201 : in_data <= 8'h9b;
      11'd1202 : in_data <= 8'h68;
      11'd1203 : in_data <= 8'hdc;
      11'd1204 : in_data <= 8'he2;
      11'd1205 : in_data <= 8'hdf;
      11'd1206 : in_data <= 8'h5e;
      11'd1207 : in_data <= 8'ha9;
      11'd1208 : in_data <= 8'h4b;
      11'd1209 : in_data <= 8'hc3;
      11'd1210 : in_data <= 8'h27;
      11'd1211 : in_data <= 8'h55;
      11'd1212 : in_data <= 8'ha5;
      11'd1213 : in_data <= 8'h97;
      11'd1214 : in_data <= 8'h66;
      11'd1215 : in_data <= 8'h4f;
      11'd1216 : in_data <= 8'hb7;
      11'd1217 : in_data <= 8'h09;
      11'd1218 : in_data <= 8'h53;
      11'd1219 : in_data <= 8'h05;
      11'd1220 : in_data <= 8'h85;
      11'd1221 : in_data <= 8'h68;
      11'd1222 : in_data <= 8'h40;
      11'd1223 : in_data <= 8'hde;
      11'd1224 : in_data <= 8'h41;
      11'd1225 : in_data <= 8'h44;
      11'd1226 : in_data <= 8'h55;
      11'd1227 : in_data <= 8'hea;
      11'd1228 : in_data <= 8'h4e;
      11'd1229 : in_data <= 8'h91;
      11'd1230 : in_data <= 8'h0a;
      11'd1231 : in_data <= 8'h21;
      11'd1232 : in_data <= 8'h34;
      11'd1233 : in_data <= 8'h86;
      11'd1234 : in_data <= 8'h40;
      11'd1235 : in_data <= 8'h8d;
      11'd1236 : in_data <= 8'h7e;
      11'd1237 : in_data <= 8'hf1;
      11'd1238 : in_data <= 8'ha3;
      11'd1239 : in_data <= 8'h6e;
      11'd1240 : in_data <= 8'h74;
      11'd1241 : in_data <= 8'h46;
      11'd1242 : in_data <= 8'hd4;
      11'd1243 : in_data <= 8'h9c;
      11'd1244 : in_data <= 8'h1d;
      11'd1245 : in_data <= 8'hd7;
      11'd1246 : in_data <= 8'ha3;
      11'd1247 : in_data <= 8'hd8;
      11'd1248 : in_data <= 8'h37;
      11'd1249 : in_data <= 8'h93;
      11'd1250 : in_data <= 8'hcc;
      11'd1251 : in_data <= 8'h2e;
      11'd1252 : in_data <= 8'he1;
      11'd1253 : in_data <= 8'h58;
      11'd1254 : in_data <= 8'h3d;
      11'd1255 : in_data <= 8'hd4;
      11'd1256 : in_data <= 8'h38;
      11'd1257 : in_data <= 8'h5f;
      11'd1258 : in_data <= 8'hd4;
      11'd1259 : in_data <= 8'h5f;
      11'd1260 : in_data <= 8'hdc;
      11'd1261 : in_data <= 8'h82;
      11'd1262 : in_data <= 8'h03;
      11'd1263 : in_data <= 8'h7b;
      11'd1264 : in_data <= 8'hd5;
      11'd1265 : in_data <= 8'h2b;
      11'd1266 : in_data <= 8'h37;
      11'd1267 : in_data <= 8'hf6;
      11'd1268 : in_data <= 8'h92;
      11'd1269 : in_data <= 8'hf8;
      11'd1270 : in_data <= 8'hc3;
      11'd1271 : in_data <= 8'h59;
      11'd1272 : in_data <= 8'hc7;
      11'd1273 : in_data <= 8'h76;
      11'd1274 : in_data <= 8'hd6;
      11'd1275 : in_data <= 8'h0e;
      11'd1276 : in_data <= 8'hf8;
      11'd1277 : in_data <= 8'h9f;
      11'd1278 : in_data <= 8'h36;
      11'd1279 : in_data <= 8'h14;
      11'd1280 : in_data <= 8'hb5;
      11'd1281 : in_data <= 8'h26;
      11'd1282 : in_data <= 8'h70;
      11'd1283 : in_data <= 8'h08;
      11'd1284 : in_data <= 8'h3a;
      11'd1285 : in_data <= 8'h06;
      11'd1286 : in_data <= 8'he7;
      11'd1287 : in_data <= 8'h39;
      11'd1288 : in_data <= 8'h3a;
      11'd1289 : in_data <= 8'h53;
      11'd1290 : in_data <= 8'h32;
      11'd1291 : in_data <= 8'hcd;
      11'd1292 : in_data <= 8'hcb;
      11'd1293 : in_data <= 8'h87;
      11'd1294 : in_data <= 8'h23;
      11'd1295 : in_data <= 8'h39;
      11'd1296 : in_data <= 8'hea;
      11'd1297 : in_data <= 8'h2b;
      11'd1298 : in_data <= 8'h35;
      11'd1299 : in_data <= 8'hd2;
      11'd1300 : in_data <= 8'hf6;
      11'd1301 : in_data <= 8'hea;
      11'd1302 : in_data <= 8'he6;
      11'd1303 : in_data <= 8'hd8;
      11'd1304 : in_data <= 8'h9a;
      11'd1305 : in_data <= 8'h03;
      11'd1306 : in_data <= 8'hc3;
      11'd1307 : in_data <= 8'h5f;
      11'd1308 : in_data <= 8'hcb;
      11'd1309 : in_data <= 8'he4;
      11'd1310 : in_data <= 8'h38;
      11'd1311 : in_data <= 8'hdd;
      11'd1312 : in_data <= 8'h9a;
      11'd1313 : in_data <= 8'hde;
      11'd1314 : in_data <= 8'h7c;
      11'd1315 : in_data <= 8'hee;
      11'd1316 : in_data <= 8'h25;
      default: in_data <= 8'h0;
    endcase
  end

  always @ ( posedge clk ) begin
    case(out_addr)
      10'd0    : out_data_ref <= 14'h0157; // 'd343
      10'd1    : out_data_ref <= 14'h00f1; // 'd241
      10'd2    : out_data_ref <= 14'h077c; // 'd1916
      10'd3    : out_data_ref <= 14'h05aa; // 'd1450
      10'd4    : out_data_ref <= 14'h0333; // 'd819
      10'd5    : out_data_ref <= 14'h0630; // 'd1584
      10'd6    : out_data_ref <= 14'h02b7; // 'd695
      10'd7    : out_data_ref <= 14'h0061; // 'd97
      10'd8    : out_data_ref <= 14'h04d0; // 'd1232
      10'd9    : out_data_ref <= 14'h0649; // 'd1609
      10'd10   : out_data_ref <= 14'h0056; // 'd86
      10'd11   : out_data_ref <= 14'h030d; // 'd781
      10'd12   : out_data_ref <= 14'h0500; // 'd1280
      10'd13   : out_data_ref <= 14'h00fc; // 'd252
      10'd14   : out_data_ref <= 14'h04d0; // 'd1232
      10'd15   : out_data_ref <= 14'h0668; // 'd1640
      10'd16   : out_data_ref <= 14'h0290; // 'd656
      10'd17   : out_data_ref <= 14'h0422; // 'd1058
      10'd18   : out_data_ref <= 14'h05bc; // 'd1468
      10'd19   : out_data_ref <= 14'h0702; // 'd1794
      10'd20   : out_data_ref <= 14'h06f7; // 'd1783
      10'd21   : out_data_ref <= 14'h04d8; // 'd1240
      10'd22   : out_data_ref <= 14'h04e4; // 'd1252
      10'd23   : out_data_ref <= 14'h07d7; // 'd2007
      10'd24   : out_data_ref <= 14'h05b3; // 'd1459
      10'd25   : out_data_ref <= 14'h0451; // 'd1105
      10'd26   : out_data_ref <= 14'h001a; // 'd26
      10'd27   : out_data_ref <= 14'h0176; // 'd374
      10'd28   : out_data_ref <= 14'h0666; // 'd1638
      10'd29   : out_data_ref <= 14'h0286; // 'd646
      10'd30   : out_data_ref <= 14'h0673; // 'd1651
      10'd31   : out_data_ref <= 14'h05ff; // 'd1535
      10'd32   : out_data_ref <= 14'h0422; // 'd1058
      10'd33   : out_data_ref <= 14'h0659; // 'd1625
      10'd34   : out_data_ref <= 14'h05df; // 'd1503
      10'd35   : out_data_ref <= 14'h0548; // 'd1352
      10'd36   : out_data_ref <= 14'h027b; // 'd635
      10'd37   : out_data_ref <= 14'h0440; // 'd1088
      10'd38   : out_data_ref <= 14'h0392; // 'd914
      10'd39   : out_data_ref <= 14'h074b; // 'd1867
      10'd40   : out_data_ref <= 14'h07ec; // 'd2028
      10'd41   : out_data_ref <= 14'h0313; // 'd787
      10'd42   : out_data_ref <= 14'h01c5; // 'd453
      10'd43   : out_data_ref <= 14'h07fc; // 'd2044
      10'd44   : out_data_ref <= 14'h054e; // 'd1358
      10'd45   : out_data_ref <= 14'h03ed; // 'd1005
      10'd46   : out_data_ref <= 14'h081c; // 'd2076
      10'd47   : out_data_ref <= 14'h008f; // 'd143
      10'd48   : out_data_ref <= 14'h0520; // 'd1312
      10'd49   : out_data_ref <= 14'h00c5; // 'd197
      10'd50   : out_data_ref <= 14'h005b; // 'd91
      10'd51   : out_data_ref <= 14'h0546; // 'd1350
      10'd52   : out_data_ref <= 14'h02d6; // 'd726
      10'd53   : out_data_ref <= 14'h053e; // 'd1342
      10'd54   : out_data_ref <= 14'h0529; // 'd1321
      10'd55   : out_data_ref <= 14'h00de; // 'd222
      10'd56   : out_data_ref <= 14'h0551; // 'd1361
      10'd57   : out_data_ref <= 14'h0388; // 'd904
      10'd58   : out_data_ref <= 14'h06c5; // 'd1733
      10'd59   : out_data_ref <= 14'h029b; // 'd667
      10'd60   : out_data_ref <= 14'h07eb; // 'd2027
      10'd61   : out_data_ref <= 14'h0246; // 'd582
      10'd62   : out_data_ref <= 14'h043f; // 'd1087
      10'd63   : out_data_ref <= 14'h045e; // 'd1118
      10'd64   : out_data_ref <= 14'h07c6; // 'd1990
      10'd65   : out_data_ref <= 14'h022c; // 'd556
      10'd66   : out_data_ref <= 14'h07c6; // 'd1990
      10'd67   : out_data_ref <= 14'h0215; // 'd533
      10'd68   : out_data_ref <= 14'h01ed; // 'd493
      10'd69   : out_data_ref <= 14'h00c2; // 'd194
      10'd70   : out_data_ref <= 14'h043b; // 'd1083
      10'd71   : out_data_ref <= 14'h0773; // 'd1907
      10'd72   : out_data_ref <= 14'h05e8; // 'd1512
      10'd73   : out_data_ref <= 14'h05dd; // 'd1501
      10'd74   : out_data_ref <= 14'h00e1; // 'd225
      10'd75   : out_data_ref <= 14'h083d; // 'd2109
      10'd76   : out_data_ref <= 14'h021c; // 'd540
      10'd77   : out_data_ref <= 14'h081d; // 'd2077
      10'd78   : out_data_ref <= 14'h01d5; // 'd469
      10'd79   : out_data_ref <= 14'h03df; // 'd991
      10'd80   : out_data_ref <= 14'h0030; // 'd48
      10'd81   : out_data_ref <= 14'h05bd; // 'd1469
      10'd82   : out_data_ref <= 14'h0520; // 'd1312
      10'd83   : out_data_ref <= 14'h05dc; // 'd1500
      10'd84   : out_data_ref <= 14'h0509; // 'd1289
      10'd85   : out_data_ref <= 14'h01a0; // 'd416
      10'd86   : out_data_ref <= 14'h0766; // 'd1894
      10'd87   : out_data_ref <= 14'h079a; // 'd1946
      10'd88   : out_data_ref <= 14'h0051; // 'd81
      10'd89   : out_data_ref <= 14'h064c; // 'd1612
      10'd90   : out_data_ref <= 14'h0180; // 'd384
      10'd91   : out_data_ref <= 14'h0657; // 'd1623
      10'd92   : out_data_ref <= 14'h0084; // 'd132
      10'd93   : out_data_ref <= 14'h03bd; // 'd957
      10'd94   : out_data_ref <= 14'h00c1; // 'd193
      10'd95   : out_data_ref <= 14'h059b; // 'd1435
      10'd96   : out_data_ref <= 14'h0331; // 'd817
      10'd97   : out_data_ref <= 14'h0418; // 'd1048
      10'd98   : out_data_ref <= 14'h066c; // 'd1644
      10'd99   : out_data_ref <= 14'h00ef; // 'd239
      10'd100  : out_data_ref <= 14'h00e6; // 'd230
      10'd101  : out_data_ref <= 14'h04c3; // 'd1219
      10'd102  : out_data_ref <= 14'h0018; // 'd24
      10'd103  : out_data_ref <= 14'h07c3; // 'd1987
      10'd104  : out_data_ref <= 14'h0645; // 'd1605
      10'd105  : out_data_ref <= 14'h070e; // 'd1806
      10'd106  : out_data_ref <= 14'h016b; // 'd363
      10'd107  : out_data_ref <= 14'h004b; // 'd75
      10'd108  : out_data_ref <= 14'h017e; // 'd382
      10'd109  : out_data_ref <= 14'h0282; // 'd642
      10'd110  : out_data_ref <= 14'h0669; // 'd1641
      10'd111  : out_data_ref <= 14'h0694; // 'd1684
      10'd112  : out_data_ref <= 14'h0636; // 'd1590
      10'd113  : out_data_ref <= 14'h0040; // 'd64
      10'd114  : out_data_ref <= 14'h0239; // 'd569
      10'd115  : out_data_ref <= 14'h03c1; // 'd961
      10'd116  : out_data_ref <= 14'h068e; // 'd1678
      10'd117  : out_data_ref <= 14'h06ea; // 'd1770
      10'd118  : out_data_ref <= 14'h0337; // 'd823
      10'd119  : out_data_ref <= 14'h00a3; // 'd163
      10'd120  : out_data_ref <= 14'h0174; // 'd372
      10'd121  : out_data_ref <= 14'h0368; // 'd872
      10'd122  : out_data_ref <= 14'h054a; // 'd1354
      10'd123  : out_data_ref <= 14'h0797; // 'd1943
      10'd124  : out_data_ref <= 14'h03ce; // 'd974
      10'd125  : out_data_ref <= 14'h0254; // 'd596
      10'd126  : out_data_ref <= 14'h07e5; // 'd2021
      10'd127  : out_data_ref <= 14'h017a; // 'd378
      10'd128  : out_data_ref <= 14'h0120; // 'd288
      10'd129  : out_data_ref <= 14'h03a5; // 'd933
      10'd130  : out_data_ref <= 14'h0210; // 'd528
      10'd131  : out_data_ref <= 14'h033b; // 'd827
      10'd132  : out_data_ref <= 14'h04bc; // 'd1212
      10'd133  : out_data_ref <= 14'h0765; // 'd1893
      10'd134  : out_data_ref <= 14'h0721; // 'd1825
      10'd135  : out_data_ref <= 14'h01d4; // 'd468
      10'd136  : out_data_ref <= 14'h0596; // 'd1430
      10'd137  : out_data_ref <= 14'h058b; // 'd1419
      10'd138  : out_data_ref <= 14'h02c2; // 'd706
      10'd139  : out_data_ref <= 14'h044f; // 'd1103
      10'd140  : out_data_ref <= 14'h0243; // 'd579
      10'd141  : out_data_ref <= 14'h046e; // 'd1134
      10'd142  : out_data_ref <= 14'h008b; // 'd139
      10'd143  : out_data_ref <= 14'h0157; // 'd343
      10'd144  : out_data_ref <= 14'h04da; // 'd1242
      10'd145  : out_data_ref <= 14'h03dc; // 'd988
      10'd146  : out_data_ref <= 14'h05e0; // 'd1504
      10'd147  : out_data_ref <= 14'h0615; // 'd1557
      10'd148  : out_data_ref <= 14'h0496; // 'd1174
      10'd149  : out_data_ref <= 14'h02d5; // 'd725
      10'd150  : out_data_ref <= 14'h04f5; // 'd1269
      10'd151  : out_data_ref <= 14'h07fb; // 'd2043
      10'd152  : out_data_ref <= 14'h0505; // 'd1285
      10'd153  : out_data_ref <= 14'h06ba; // 'd1722
      10'd154  : out_data_ref <= 14'h03f0; // 'd1008
      10'd155  : out_data_ref <= 14'h0419; // 'd1049
      10'd156  : out_data_ref <= 14'h02d6; // 'd726
      10'd157  : out_data_ref <= 14'h0600; // 'd1536
      10'd158  : out_data_ref <= 14'h05ec; // 'd1516
      10'd159  : out_data_ref <= 14'h0272; // 'd626
      10'd160  : out_data_ref <= 14'h079c; // 'd1948
      10'd161  : out_data_ref <= 14'h01d9; // 'd473
      10'd162  : out_data_ref <= 14'h0730; // 'd1840
      10'd163  : out_data_ref <= 14'h0735; // 'd1845
      10'd164  : out_data_ref <= 14'h067f; // 'd1663
      10'd165  : out_data_ref <= 14'h0544; // 'd1348
      10'd166  : out_data_ref <= 14'h06ac; // 'd1708
      10'd167  : out_data_ref <= 14'h07cf; // 'd1999
      10'd168  : out_data_ref <= 14'h002f; // 'd47
      10'd169  : out_data_ref <= 14'h002d; // 'd45
      10'd170  : out_data_ref <= 14'h021f; // 'd543
      10'd171  : out_data_ref <= 14'h0717; // 'd1815
      10'd172  : out_data_ref <= 14'h037f; // 'd895
      10'd173  : out_data_ref <= 14'h0684; // 'd1668
      10'd174  : out_data_ref <= 14'h038f; // 'd911
      10'd175  : out_data_ref <= 14'h0424; // 'd1060
      10'd176  : out_data_ref <= 14'h0082; // 'd130
      10'd177  : out_data_ref <= 14'h01fa; // 'd506
      10'd178  : out_data_ref <= 14'h0565; // 'd1381
      10'd179  : out_data_ref <= 14'h0300; // 'd768
      10'd180  : out_data_ref <= 14'h00e4; // 'd228
      10'd181  : out_data_ref <= 14'h0531; // 'd1329
      10'd182  : out_data_ref <= 14'h0558; // 'd1368
      10'd183  : out_data_ref <= 14'h0475; // 'd1141
      10'd184  : out_data_ref <= 14'h0770; // 'd1904
      10'd185  : out_data_ref <= 14'h053b; // 'd1339
      10'd186  : out_data_ref <= 14'h0180; // 'd384
      10'd187  : out_data_ref <= 14'h0537; // 'd1335
      10'd188  : out_data_ref <= 14'h0668; // 'd1640
      10'd189  : out_data_ref <= 14'h000d; // 'd13
      10'd190  : out_data_ref <= 14'h0817; // 'd2071
      10'd191  : out_data_ref <= 14'h0617; // 'd1559
      10'd192  : out_data_ref <= 14'h029a; // 'd666
      10'd193  : out_data_ref <= 14'h00ae; // 'd174
      10'd194  : out_data_ref <= 14'h0287; // 'd647
      10'd195  : out_data_ref <= 14'h0121; // 'd289
      10'd196  : out_data_ref <= 14'h00c3; // 'd195
      10'd197  : out_data_ref <= 14'h06ac; // 'd1708
      10'd198  : out_data_ref <= 14'h0768; // 'd1896
      10'd199  : out_data_ref <= 14'h070f; // 'd1807
      10'd200  : out_data_ref <= 14'h0608; // 'd1544
      10'd201  : out_data_ref <= 14'h05e2; // 'd1506
      10'd202  : out_data_ref <= 14'h028e; // 'd654
      10'd203  : out_data_ref <= 14'h082d; // 'd2093
      10'd204  : out_data_ref <= 14'h0694; // 'd1684
      10'd205  : out_data_ref <= 14'h07ed; // 'd2029
      10'd206  : out_data_ref <= 14'h01af; // 'd431
      10'd207  : out_data_ref <= 14'h07c0; // 'd1984
      10'd208  : out_data_ref <= 14'h022e; // 'd558
      10'd209  : out_data_ref <= 14'h0164; // 'd356
      10'd210  : out_data_ref <= 14'h0359; // 'd857
      10'd211  : out_data_ref <= 14'h0577; // 'd1399
      10'd212  : out_data_ref <= 14'h033c; // 'd828
      10'd213  : out_data_ref <= 14'h07d6; // 'd2006
      10'd214  : out_data_ref <= 14'h07f8; // 'd2040
      10'd215  : out_data_ref <= 14'h060c; // 'd1548
      10'd216  : out_data_ref <= 14'h04f0; // 'd1264
      10'd217  : out_data_ref <= 14'h06d1; // 'd1745
      10'd218  : out_data_ref <= 14'h0619; // 'd1561
      10'd219  : out_data_ref <= 14'h06f4; // 'd1780
      10'd220  : out_data_ref <= 14'h07e0; // 'd2016
      10'd221  : out_data_ref <= 14'h0477; // 'd1143
      10'd222  : out_data_ref <= 14'h083b; // 'd2107
      10'd223  : out_data_ref <= 14'h0530; // 'd1328
      10'd224  : out_data_ref <= 14'h0324; // 'd804
      10'd225  : out_data_ref <= 14'h0028; // 'd40
      10'd226  : out_data_ref <= 14'h02c3; // 'd707
      10'd227  : out_data_ref <= 14'h0570; // 'd1392
      10'd228  : out_data_ref <= 14'h0072; // 'd114
      10'd229  : out_data_ref <= 14'h0613; // 'd1555
      10'd230  : out_data_ref <= 14'h017b; // 'd379
      10'd231  : out_data_ref <= 14'h0755; // 'd1877
      10'd232  : out_data_ref <= 14'h0839; // 'd2105
      10'd233  : out_data_ref <= 14'h07cd; // 'd1997
      10'd234  : out_data_ref <= 14'h07fa; // 'd2042
      10'd235  : out_data_ref <= 14'h049f; // 'd1183
      10'd236  : out_data_ref <= 14'h04be; // 'd1214
      10'd237  : out_data_ref <= 14'h0175; // 'd373
      10'd238  : out_data_ref <= 14'h0516; // 'd1302
      10'd239  : out_data_ref <= 14'h055c; // 'd1372
      10'd240  : out_data_ref <= 14'h01a7; // 'd423
      10'd241  : out_data_ref <= 14'h0836; // 'd2102
      10'd242  : out_data_ref <= 14'h0744; // 'd1860
      10'd243  : out_data_ref <= 14'h053e; // 'd1342
      10'd244  : out_data_ref <= 14'h01a3; // 'd419
      10'd245  : out_data_ref <= 14'h0676; // 'd1654
      10'd246  : out_data_ref <= 14'h06ae; // 'd1710
      10'd247  : out_data_ref <= 14'h01e7; // 'd487
      10'd248  : out_data_ref <= 14'h0671; // 'd1649
      10'd249  : out_data_ref <= 14'h05e9; // 'd1513
      10'd250  : out_data_ref <= 14'h04c7; // 'd1223
      10'd251  : out_data_ref <= 14'h067f; // 'd1663
      10'd252  : out_data_ref <= 14'h055e; // 'd1374
      10'd253  : out_data_ref <= 14'h0369; // 'd873
      10'd254  : out_data_ref <= 14'h083c; // 'd2108
      10'd255  : out_data_ref <= 14'h0598; // 'd1432
      10'd256  : out_data_ref <= 14'h062c; // 'd1580
      10'd257  : out_data_ref <= 14'h082c; // 'd2092
      10'd258  : out_data_ref <= 14'h06d2; // 'd1746
      10'd259  : out_data_ref <= 14'h00e5; // 'd229
      10'd260  : out_data_ref <= 14'h0399; // 'd921
      10'd261  : out_data_ref <= 14'h0297; // 'd663
      10'd262  : out_data_ref <= 14'h077b; // 'd1915
      10'd263  : out_data_ref <= 14'h01e7; // 'd487
      10'd264  : out_data_ref <= 14'h006b; // 'd107
      10'd265  : out_data_ref <= 14'h05db; // 'd1499
      10'd266  : out_data_ref <= 14'h0609; // 'd1545
      10'd267  : out_data_ref <= 14'h04c7; // 'd1223
      10'd268  : out_data_ref <= 14'h03f7; // 'd1015
      10'd269  : out_data_ref <= 14'h0459; // 'd1113
      10'd270  : out_data_ref <= 14'h01de; // 'd478
      10'd271  : out_data_ref <= 14'h01d9; // 'd473
      10'd272  : out_data_ref <= 14'h000c; // 'd12
      10'd273  : out_data_ref <= 14'h04ba; // 'd1210
      10'd274  : out_data_ref <= 14'h00c5; // 'd197
      10'd275  : out_data_ref <= 14'h0747; // 'd1863
      10'd276  : out_data_ref <= 14'h0082; // 'd130
      10'd277  : out_data_ref <= 14'h04a2; // 'd1186
      10'd278  : out_data_ref <= 14'h0414; // 'd1044
      10'd279  : out_data_ref <= 14'h055a; // 'd1370
      10'd280  : out_data_ref <= 14'h075f; // 'd1887
      10'd281  : out_data_ref <= 14'h03ca; // 'd970
      10'd282  : out_data_ref <= 14'h039a; // 'd922
      10'd283  : out_data_ref <= 14'h00b0; // 'd176
      10'd284  : out_data_ref <= 14'h00a7; // 'd167
      10'd285  : out_data_ref <= 14'h04ed; // 'd1261
      10'd286  : out_data_ref <= 14'h0298; // 'd664
      10'd287  : out_data_ref <= 14'h03bc; // 'd956
      10'd288  : out_data_ref <= 14'h0057; // 'd87
      10'd289  : out_data_ref <= 14'h053a; // 'd1338
      10'd290  : out_data_ref <= 14'h07b4; // 'd1972
      10'd291  : out_data_ref <= 14'h0764; // 'd1892
      10'd292  : out_data_ref <= 14'h0324; // 'd804
      10'd293  : out_data_ref <= 14'h015d; // 'd349
      10'd294  : out_data_ref <= 14'h031d; // 'd797
      10'd295  : out_data_ref <= 14'h0752; // 'd1874
      10'd296  : out_data_ref <= 14'h0560; // 'd1376
      10'd297  : out_data_ref <= 14'h0167; // 'd359
      10'd298  : out_data_ref <= 14'h02af; // 'd687
      10'd299  : out_data_ref <= 14'h058a; // 'd1418
      10'd300  : out_data_ref <= 14'h06ea; // 'd1770
      10'd301  : out_data_ref <= 14'h067f; // 'd1663
      10'd302  : out_data_ref <= 14'h04c6; // 'd1222
      10'd303  : out_data_ref <= 14'h0101; // 'd257
      10'd304  : out_data_ref <= 14'h036f; // 'd879
      10'd305  : out_data_ref <= 14'h028e; // 'd654
      10'd306  : out_data_ref <= 14'h006a; // 'd106
      10'd307  : out_data_ref <= 14'h0197; // 'd407
      10'd308  : out_data_ref <= 14'h030e; // 'd782
      10'd309  : out_data_ref <= 14'h01c6; // 'd454
      10'd310  : out_data_ref <= 14'h0152; // 'd338
      10'd311  : out_data_ref <= 14'h02ae; // 'd686
      10'd312  : out_data_ref <= 14'h05a1; // 'd1441
      10'd313  : out_data_ref <= 14'h07bd; // 'd1981
      10'd314  : out_data_ref <= 14'h0265; // 'd613
      10'd315  : out_data_ref <= 14'h055d; // 'd1373
      10'd316  : out_data_ref <= 14'h0047; // 'd71
      10'd317  : out_data_ref <= 14'h0218; // 'd536
      10'd318  : out_data_ref <= 14'h07d2; // 'd2002
      10'd319  : out_data_ref <= 14'h0385; // 'd901
      10'd320  : out_data_ref <= 14'h00fb; // 'd251
      10'd321  : out_data_ref <= 14'h03f6; // 'd1014
      10'd322  : out_data_ref <= 14'h0460; // 'd1120
      10'd323  : out_data_ref <= 14'h027e; // 'd638
      10'd324  : out_data_ref <= 14'h0078; // 'd120
      10'd325  : out_data_ref <= 14'h033e; // 'd830
      10'd326  : out_data_ref <= 14'h00a1; // 'd161
      10'd327  : out_data_ref <= 14'h077a; // 'd1914
      10'd328  : out_data_ref <= 14'h06fe; // 'd1790
      10'd329  : out_data_ref <= 14'h05d1; // 'd1489
      10'd330  : out_data_ref <= 14'h0032; // 'd50
      10'd331  : out_data_ref <= 14'h04de; // 'd1246
      10'd332  : out_data_ref <= 14'h033c; // 'd828
      10'd333  : out_data_ref <= 14'h03bc; // 'd956
      10'd334  : out_data_ref <= 14'h0622; // 'd1570
      10'd335  : out_data_ref <= 14'h03ea; // 'd1002
      10'd336  : out_data_ref <= 14'h003d; // 'd61
      10'd337  : out_data_ref <= 14'h00d3; // 'd211
      10'd338  : out_data_ref <= 14'h078f; // 'd1935
      10'd339  : out_data_ref <= 14'h0616; // 'd1558
      10'd340  : out_data_ref <= 14'h053f; // 'd1343
      10'd341  : out_data_ref <= 14'h0001; // 'd1
      10'd342  : out_data_ref <= 14'h06bb; // 'd1723
      10'd343  : out_data_ref <= 14'h031b; // 'd795
      10'd344  : out_data_ref <= 14'h0650; // 'd1616
      10'd345  : out_data_ref <= 14'h00e9; // 'd233
      10'd346  : out_data_ref <= 14'h0793; // 'd1939
      10'd347  : out_data_ref <= 14'h082c; // 'd2092
      10'd348  : out_data_ref <= 14'h04fb; // 'd1275
      10'd349  : out_data_ref <= 14'h0664; // 'd1636
      10'd350  : out_data_ref <= 14'h06d6; // 'd1750
      10'd351  : out_data_ref <= 14'h06c7; // 'd1735
      10'd352  : out_data_ref <= 14'h058f; // 'd1423
      10'd353  : out_data_ref <= 14'h02fe; // 'd766
      10'd354  : out_data_ref <= 14'h0634; // 'd1588
      10'd355  : out_data_ref <= 14'h05b3; // 'd1459
      10'd356  : out_data_ref <= 14'h041c; // 'd1052
      10'd357  : out_data_ref <= 14'h03a8; // 'd936
      10'd358  : out_data_ref <= 14'h0441; // 'd1089
      10'd359  : out_data_ref <= 14'h0297; // 'd663
      10'd360  : out_data_ref <= 14'h077d; // 'd1917
      10'd361  : out_data_ref <= 14'h00ee; // 'd238
      10'd362  : out_data_ref <= 14'h04a8; // 'd1192
      10'd363  : out_data_ref <= 14'h0079; // 'd121
      10'd364  : out_data_ref <= 14'h02ac; // 'd684
      10'd365  : out_data_ref <= 14'h073b; // 'd1851
      10'd366  : out_data_ref <= 14'h049e; // 'd1182
      10'd367  : out_data_ref <= 14'h0121; // 'd289
      10'd368  : out_data_ref <= 14'h01e8; // 'd488
      10'd369  : out_data_ref <= 14'h07a0; // 'd1952
      10'd370  : out_data_ref <= 14'h00b1; // 'd177
      10'd371  : out_data_ref <= 14'h07e8; // 'd2024
      10'd372  : out_data_ref <= 14'h0683; // 'd1667
      10'd373  : out_data_ref <= 14'h0802; // 'd2050
      10'd374  : out_data_ref <= 14'h03af; // 'd943
      10'd375  : out_data_ref <= 14'h032b; // 'd811
      10'd376  : out_data_ref <= 14'h06a0; // 'd1696
      10'd377  : out_data_ref <= 14'h027f; // 'd639
      10'd378  : out_data_ref <= 14'h04d4; // 'd1236
      10'd379  : out_data_ref <= 14'h0718; // 'd1816
      10'd380  : out_data_ref <= 14'h0064; // 'd100
      10'd381  : out_data_ref <= 14'h0091; // 'd145
      10'd382  : out_data_ref <= 14'h030d; // 'd781
      10'd383  : out_data_ref <= 14'h0736; // 'd1846
      10'd384  : out_data_ref <= 14'h0131; // 'd305
      10'd385  : out_data_ref <= 14'h06db; // 'd1755
      10'd386  : out_data_ref <= 14'h0323; // 'd803
      10'd387  : out_data_ref <= 14'h06b8; // 'd1720
      10'd388  : out_data_ref <= 14'h019e; // 'd414
      10'd389  : out_data_ref <= 14'h0568; // 'd1384
      10'd390  : out_data_ref <= 14'h03e2; // 'd994
      10'd391  : out_data_ref <= 14'h0386; // 'd902
      10'd392  : out_data_ref <= 14'h0484; // 'd1156
      10'd393  : out_data_ref <= 14'h033d; // 'd829
      10'd394  : out_data_ref <= 14'h0294; // 'd660
      10'd395  : out_data_ref <= 14'h0800; // 'd2048
      10'd396  : out_data_ref <= 14'h03cd; // 'd973
      10'd397  : out_data_ref <= 14'h0062; // 'd98
      10'd398  : out_data_ref <= 14'h081f; // 'd2079
      10'd399  : out_data_ref <= 14'h0749; // 'd1865
      10'd400  : out_data_ref <= 14'h01e4; // 'd484
      10'd401  : out_data_ref <= 14'h0382; // 'd898
      10'd402  : out_data_ref <= 14'h02e6; // 'd742
      10'd403  : out_data_ref <= 14'h0373; // 'd883
      10'd404  : out_data_ref <= 14'h049f; // 'd1183
      10'd405  : out_data_ref <= 14'h01d1; // 'd465
      10'd406  : out_data_ref <= 14'h0684; // 'd1668
      10'd407  : out_data_ref <= 14'h0057; // 'd87
      10'd408  : out_data_ref <= 14'h05d9; // 'd1497
      10'd409  : out_data_ref <= 14'h016a; // 'd362
      10'd410  : out_data_ref <= 14'h0558; // 'd1368
      10'd411  : out_data_ref <= 14'h0051; // 'd81
      10'd412  : out_data_ref <= 14'h00d3; // 'd211
      10'd413  : out_data_ref <= 14'h01d9; // 'd473
      10'd414  : out_data_ref <= 14'h00ef; // 'd239
      10'd415  : out_data_ref <= 14'h02a0; // 'd672
      10'd416  : out_data_ref <= 14'h07c1; // 'd1985
      10'd417  : out_data_ref <= 14'h01d9; // 'd473
      10'd418  : out_data_ref <= 14'h0243; // 'd579
      10'd419  : out_data_ref <= 14'h0506; // 'd1286
      10'd420  : out_data_ref <= 14'h03d9; // 'd985
      10'd421  : out_data_ref <= 14'h027c; // 'd636
      10'd422  : out_data_ref <= 14'h0628; // 'd1576
      10'd423  : out_data_ref <= 14'h0144; // 'd324
      10'd424  : out_data_ref <= 14'h02a9; // 'd681
      10'd425  : out_data_ref <= 14'h04f4; // 'd1268
      10'd426  : out_data_ref <= 14'h0668; // 'd1640
      10'd427  : out_data_ref <= 14'h04b2; // 'd1202
      10'd428  : out_data_ref <= 14'h059f; // 'd1439
      10'd429  : out_data_ref <= 14'h0202; // 'd514
      10'd430  : out_data_ref <= 14'h0261; // 'd609
      10'd431  : out_data_ref <= 14'h0673; // 'd1651
      10'd432  : out_data_ref <= 14'h035a; // 'd858
      10'd433  : out_data_ref <= 14'h03bf; // 'd959
      10'd434  : out_data_ref <= 14'h00ee; // 'd238
      10'd435  : out_data_ref <= 14'h079f; // 'd1951
      10'd436  : out_data_ref <= 14'h05d6; // 'd1494
      10'd437  : out_data_ref <= 14'h0051; // 'd81
      10'd438  : out_data_ref <= 14'h0060; // 'd96
      10'd439  : out_data_ref <= 14'h002d; // 'd45
      10'd440  : out_data_ref <= 14'h0608; // 'd1544
      10'd441  : out_data_ref <= 14'h0223; // 'd547
      10'd442  : out_data_ref <= 14'h06a9; // 'd1705
      10'd443  : out_data_ref <= 14'h05ca; // 'd1482
      10'd444  : out_data_ref <= 14'h0776; // 'd1910
      10'd445  : out_data_ref <= 14'h039f; // 'd927
      10'd446  : out_data_ref <= 14'h0130; // 'd304
      10'd447  : out_data_ref <= 14'h04db; // 'd1243
      10'd448  : out_data_ref <= 14'h00dc; // 'd220
      10'd449  : out_data_ref <= 14'h0734; // 'd1844
      10'd450  : out_data_ref <= 14'h05a4; // 'd1444
      10'd451  : out_data_ref <= 14'h0530; // 'd1328
      10'd452  : out_data_ref <= 14'h01d0; // 'd464
      10'd453  : out_data_ref <= 14'h02d1; // 'd721
      10'd454  : out_data_ref <= 14'h072d; // 'd1837
      10'd455  : out_data_ref <= 14'h05fb; // 'd1531
      10'd456  : out_data_ref <= 14'h03d5; // 'd981
      10'd457  : out_data_ref <= 14'h064f; // 'd1615
      10'd458  : out_data_ref <= 14'h05ba; // 'd1466
      10'd459  : out_data_ref <= 14'h01be; // 'd446
      10'd460  : out_data_ref <= 14'h072f; // 'd1839
      10'd461  : out_data_ref <= 14'h012e; // 'd302
      10'd462  : out_data_ref <= 14'h0169; // 'd361
      10'd463  : out_data_ref <= 14'h041d; // 'd1053
      10'd464  : out_data_ref <= 14'h0001; // 'd1
      10'd465  : out_data_ref <= 14'h0689; // 'd1673
      10'd466  : out_data_ref <= 14'h063d; // 'd1597
      10'd467  : out_data_ref <= 14'h0338; // 'd824
      10'd468  : out_data_ref <= 14'h0177; // 'd375
      10'd469  : out_data_ref <= 14'h0146; // 'd326
      10'd470  : out_data_ref <= 14'h054c; // 'd1356
      10'd471  : out_data_ref <= 14'h03f0; // 'd1008
      10'd472  : out_data_ref <= 14'h0826; // 'd2086
      10'd473  : out_data_ref <= 14'h00f8; // 'd248
      10'd474  : out_data_ref <= 14'h0721; // 'd1825
      10'd475  : out_data_ref <= 14'h04d3; // 'd1235
      10'd476  : out_data_ref <= 14'h0817; // 'd2071
      10'd477  : out_data_ref <= 14'h05f2; // 'd1522
      10'd478  : out_data_ref <= 14'h04d4; // 'd1236
      10'd479  : out_data_ref <= 14'h0795; // 'd1941
      10'd480  : out_data_ref <= 14'h00a2; // 'd162
      10'd481  : out_data_ref <= 14'h0002; // 'd2
      10'd482  : out_data_ref <= 14'h0721; // 'd1825
      10'd483  : out_data_ref <= 14'h0613; // 'd1555
      10'd484  : out_data_ref <= 14'h0558; // 'd1368
      10'd485  : out_data_ref <= 14'h025e; // 'd606
      10'd486  : out_data_ref <= 14'h0587; // 'd1415
      10'd487  : out_data_ref <= 14'h0333; // 'd819
      10'd488  : out_data_ref <= 14'h02e6; // 'd742
      10'd489  : out_data_ref <= 14'h01db; // 'd475
      10'd490  : out_data_ref <= 14'h05c2; // 'd1474
      10'd491  : out_data_ref <= 14'h0749; // 'd1865
      10'd492  : out_data_ref <= 14'h0288; // 'd648
      10'd493  : out_data_ref <= 14'h00a6; // 'd166
      10'd494  : out_data_ref <= 14'h03dc; // 'd988
      10'd495  : out_data_ref <= 14'h040b; // 'd1035
      10'd496  : out_data_ref <= 14'h047c; // 'd1148
      10'd497  : out_data_ref <= 14'h066b; // 'd1643
      10'd498  : out_data_ref <= 14'h062f; // 'd1583
      10'd499  : out_data_ref <= 14'h0646; // 'd1606
      10'd500  : out_data_ref <= 14'h03ac; // 'd940
      10'd501  : out_data_ref <= 14'h0526; // 'd1318
      10'd502  : out_data_ref <= 14'h021c; // 'd540
      10'd503  : out_data_ref <= 14'h072e; // 'd1838
      10'd504  : out_data_ref <= 14'h051f; // 'd1311
      10'd505  : out_data_ref <= 14'h077f; // 'd1919
      10'd506  : out_data_ref <= 14'h00d5; // 'd213
      10'd507  : out_data_ref <= 14'h06d6; // 'd1750
      10'd508  : out_data_ref <= 14'h0075; // 'd117
      10'd509  : out_data_ref <= 14'h04fb; // 'd1275
      10'd510  : out_data_ref <= 14'h00ac; // 'd172
      10'd511  : out_data_ref <= 14'h0305; // 'd773
      10'd512  : out_data_ref <= 14'h052d; // 'd1325
      10'd513  : out_data_ref <= 14'h07bd; // 'd1981
      10'd514  : out_data_ref <= 14'h045b; // 'd1115
      10'd515  : out_data_ref <= 14'h006a; // 'd106
      10'd516  : out_data_ref <= 14'h048e; // 'd1166
      10'd517  : out_data_ref <= 14'h05a2; // 'd1442
      10'd518  : out_data_ref <= 14'h0404; // 'd1028
      10'd519  : out_data_ref <= 14'h026b; // 'd619
      10'd520  : out_data_ref <= 14'h00f7; // 'd247
      10'd521  : out_data_ref <= 14'h0520; // 'd1312
      10'd522  : out_data_ref <= 14'h055e; // 'd1374
      10'd523  : out_data_ref <= 14'h0175; // 'd373
      10'd524  : out_data_ref <= 14'h052f; // 'd1327
      10'd525  : out_data_ref <= 14'h0343; // 'd835
      10'd526  : out_data_ref <= 14'h0545; // 'd1349
      10'd527  : out_data_ref <= 14'h0052; // 'd82
      10'd528  : out_data_ref <= 14'h0619; // 'd1561
      10'd529  : out_data_ref <= 14'h01df; // 'd479
      10'd530  : out_data_ref <= 14'h033d; // 'd829
      10'd531  : out_data_ref <= 14'h0429; // 'd1065
      10'd532  : out_data_ref <= 14'h059b; // 'd1435
      10'd533  : out_data_ref <= 14'h04a9; // 'd1193
      10'd534  : out_data_ref <= 14'h017f; // 'd383
      10'd535  : out_data_ref <= 14'h01ce; // 'd462
      10'd536  : out_data_ref <= 14'h0780; // 'd1920
      10'd537  : out_data_ref <= 14'h03a5; // 'd933
      10'd538  : out_data_ref <= 14'h0510; // 'd1296
      10'd539  : out_data_ref <= 14'h0100; // 'd256
      10'd540  : out_data_ref <= 14'h010b; // 'd267
      10'd541  : out_data_ref <= 14'h083d; // 'd2109
      10'd542  : out_data_ref <= 14'h054b; // 'd1355
      10'd543  : out_data_ref <= 14'h052d; // 'd1325
      10'd544  : out_data_ref <= 14'h06f4; // 'd1780
      10'd545  : out_data_ref <= 14'h0520; // 'd1312
      10'd546  : out_data_ref <= 14'h04ae; // 'd1198
      10'd547  : out_data_ref <= 14'h080d; // 'd2061
      10'd548  : out_data_ref <= 14'h07eb; // 'd2027
      10'd549  : out_data_ref <= 14'h01ad; // 'd429
      10'd550  : out_data_ref <= 14'h01ff; // 'd511
      10'd551  : out_data_ref <= 14'h0141; // 'd321
      10'd552  : out_data_ref <= 14'h056d; // 'd1389
      10'd553  : out_data_ref <= 14'h04ce; // 'd1230
      10'd554  : out_data_ref <= 14'h023b; // 'd571
      10'd555  : out_data_ref <= 14'h03c9; // 'd969
      10'd556  : out_data_ref <= 14'h0442; // 'd1090
      10'd557  : out_data_ref <= 14'h05cf; // 'd1487
      10'd558  : out_data_ref <= 14'h059e; // 'd1438
      10'd559  : out_data_ref <= 14'h062f; // 'd1583
      10'd560  : out_data_ref <= 14'h0364; // 'd868
      10'd561  : out_data_ref <= 14'h00cf; // 'd207
      10'd562  : out_data_ref <= 14'h014e; // 'd334
      10'd563  : out_data_ref <= 14'h031a; // 'd794
      10'd564  : out_data_ref <= 14'h0018; // 'd24
      10'd565  : out_data_ref <= 14'h05d5; // 'd1493
      10'd566  : out_data_ref <= 14'h0215; // 'd533
      10'd567  : out_data_ref <= 14'h0796; // 'd1942
      10'd568  : out_data_ref <= 14'h0384; // 'd900
      10'd569  : out_data_ref <= 14'h0316; // 'd790
      10'd570  : out_data_ref <= 14'h06fa; // 'd1786
      10'd571  : out_data_ref <= 14'h0384; // 'd900
      10'd572  : out_data_ref <= 14'h05aa; // 'd1450
      10'd573  : out_data_ref <= 14'h0438; // 'd1080
      10'd574  : out_data_ref <= 14'h03c5; // 'd965
      10'd575  : out_data_ref <= 14'h0168; // 'd360
      10'd576  : out_data_ref <= 14'h0138; // 'd312
      10'd577  : out_data_ref <= 14'h01aa; // 'd426
      10'd578  : out_data_ref <= 14'h05e4; // 'd1508
      10'd579  : out_data_ref <= 14'h019d; // 'd413
      10'd580  : out_data_ref <= 14'h02b5; // 'd693
      10'd581  : out_data_ref <= 14'h066c; // 'd1644
      10'd582  : out_data_ref <= 14'h05cf; // 'd1487
      10'd583  : out_data_ref <= 14'h0542; // 'd1346
      10'd584  : out_data_ref <= 14'h0155; // 'd341
      10'd585  : out_data_ref <= 14'h05b7; // 'd1463
      10'd586  : out_data_ref <= 14'h053b; // 'd1339
      10'd587  : out_data_ref <= 14'h02c0; // 'd704
      10'd588  : out_data_ref <= 14'h075f; // 'd1887
      10'd589  : out_data_ref <= 14'h026d; // 'd621
      10'd590  : out_data_ref <= 14'h052c; // 'd1324
      10'd591  : out_data_ref <= 14'h01fa; // 'd506
      10'd592  : out_data_ref <= 14'h0704; // 'd1796
      10'd593  : out_data_ref <= 14'h0544; // 'd1348
      10'd594  : out_data_ref <= 14'h0172; // 'd370
      10'd595  : out_data_ref <= 14'h0760; // 'd1888
      10'd596  : out_data_ref <= 14'h00e3; // 'd227
      10'd597  : out_data_ref <= 14'h05ce; // 'd1486
      10'd598  : out_data_ref <= 14'h0761; // 'd1889
      10'd599  : out_data_ref <= 14'h00af; // 'd175
      10'd600  : out_data_ref <= 14'h013e; // 'd318
      10'd601  : out_data_ref <= 14'h003e; // 'd62
      10'd602  : out_data_ref <= 14'h0576; // 'd1398
      10'd603  : out_data_ref <= 14'h07c7; // 'd1991
      10'd604  : out_data_ref <= 14'h07d1; // 'd2001
      10'd605  : out_data_ref <= 14'h0661; // 'd1633
      10'd606  : out_data_ref <= 14'h047c; // 'd1148
      10'd607  : out_data_ref <= 14'h0263; // 'd611
      10'd608  : out_data_ref <= 14'h0239; // 'd569
      10'd609  : out_data_ref <= 14'h00cc; // 'd204
      10'd610  : out_data_ref <= 14'h07e2; // 'd2018
      10'd611  : out_data_ref <= 14'h021b; // 'd539
      10'd612  : out_data_ref <= 14'h0507; // 'd1287
      10'd613  : out_data_ref <= 14'h00ab; // 'd171
      10'd614  : out_data_ref <= 14'h0731; // 'd1841
      10'd615  : out_data_ref <= 14'h05a7; // 'd1447
      10'd616  : out_data_ref <= 14'h04cf; // 'd1231
      10'd617  : out_data_ref <= 14'h0040; // 'd64
      10'd618  : out_data_ref <= 14'h076e; // 'd1902
      10'd619  : out_data_ref <= 14'h07ab; // 'd1963
      10'd620  : out_data_ref <= 14'h0083; // 'd131
      10'd621  : out_data_ref <= 14'h0065; // 'd101
      10'd622  : out_data_ref <= 14'h0702; // 'd1794
      10'd623  : out_data_ref <= 14'h0651; // 'd1617
      10'd624  : out_data_ref <= 14'h0430; // 'd1072
      10'd625  : out_data_ref <= 14'h0377; // 'd887
      10'd626  : out_data_ref <= 14'h03fd; // 'd1021
      10'd627  : out_data_ref <= 14'h03a7; // 'd935
      10'd628  : out_data_ref <= 14'h0312; // 'd786
      10'd629  : out_data_ref <= 14'h02c3; // 'd707
      10'd630  : out_data_ref <= 14'h03eb; // 'd1003
      10'd631  : out_data_ref <= 14'h0409; // 'd1033
      10'd632  : out_data_ref <= 14'h02af; // 'd687
      10'd633  : out_data_ref <= 14'h0553; // 'd1363
      10'd634  : out_data_ref <= 14'h0046; // 'd70
      10'd635  : out_data_ref <= 14'h0449; // 'd1097
      10'd636  : out_data_ref <= 14'h038a; // 'd906
      10'd637  : out_data_ref <= 14'h07f2; // 'd2034
      10'd638  : out_data_ref <= 14'h0109; // 'd265
      10'd639  : out_data_ref <= 14'h0275; // 'd629
      10'd640  : out_data_ref <= 14'h0712; // 'd1810
      10'd641  : out_data_ref <= 14'h06e3; // 'd1763
      10'd642  : out_data_ref <= 14'h04a1; // 'd1185
      10'd643  : out_data_ref <= 14'h0241; // 'd577
      10'd644  : out_data_ref <= 14'h030a; // 'd778
      10'd645  : out_data_ref <= 14'h06b0; // 'd1712
      10'd646  : out_data_ref <= 14'h0059; // 'd89
      10'd647  : out_data_ref <= 14'h083e; // 'd2110
      10'd648  : out_data_ref <= 14'h036a; // 'd874
      10'd649  : out_data_ref <= 14'h05ab; // 'd1451
      10'd650  : out_data_ref <= 14'h02e8; // 'd744
      10'd651  : out_data_ref <= 14'h0384; // 'd900
      10'd652  : out_data_ref <= 14'h0464; // 'd1124
      10'd653  : out_data_ref <= 14'h05ed; // 'd1517
      10'd654  : out_data_ref <= 14'h06df; // 'd1759
      10'd655  : out_data_ref <= 14'h024a; // 'd586
      10'd656  : out_data_ref <= 14'h0426; // 'd1062
      10'd657  : out_data_ref <= 14'h0681; // 'd1665
      10'd658  : out_data_ref <= 14'h043e; // 'd1086
      10'd659  : out_data_ref <= 14'h0314; // 'd788
      10'd660  : out_data_ref <= 14'h0495; // 'd1173
      10'd661  : out_data_ref <= 14'h0003; // 'd3
      10'd662  : out_data_ref <= 14'h05cb; // 'd1483
      10'd663  : out_data_ref <= 14'h0360; // 'd864
      10'd664  : out_data_ref <= 14'h043a; // 'd1082
      10'd665  : out_data_ref <= 14'h07c8; // 'd1992
      10'd666  : out_data_ref <= 14'h0372; // 'd882
      10'd667  : out_data_ref <= 14'h0394; // 'd916
      10'd668  : out_data_ref <= 14'h0675; // 'd1653
      10'd669  : out_data_ref <= 14'h066d; // 'd1645
      10'd670  : out_data_ref <= 14'h0426; // 'd1062
      10'd671  : out_data_ref <= 14'h00c1; // 'd193
      10'd672  : out_data_ref <= 14'h0287; // 'd647
      10'd673  : out_data_ref <= 14'h0421; // 'd1057
      10'd674  : out_data_ref <= 14'h06c9; // 'd1737
      10'd675  : out_data_ref <= 14'h007a; // 'd122
      10'd676  : out_data_ref <= 14'h03e3; // 'd995
      10'd677  : out_data_ref <= 14'h0047; // 'd71
      10'd678  : out_data_ref <= 14'h0296; // 'd662
      10'd679  : out_data_ref <= 14'h071e; // 'd1822
      10'd680  : out_data_ref <= 14'h045d; // 'd1117
      10'd681  : out_data_ref <= 14'h0757; // 'd1879
      10'd682  : out_data_ref <= 14'h0138; // 'd312
      10'd683  : out_data_ref <= 14'h02a0; // 'd672
      10'd684  : out_data_ref <= 14'h01bb; // 'd443
      10'd685  : out_data_ref <= 14'h0353; // 'd851
      10'd686  : out_data_ref <= 14'h04b3; // 'd1203
      10'd687  : out_data_ref <= 14'h01ef; // 'd495
      10'd688  : out_data_ref <= 14'h077f; // 'd1919
      10'd689  : out_data_ref <= 14'h0723; // 'd1827
      10'd690  : out_data_ref <= 14'h05ba; // 'd1466
      10'd691  : out_data_ref <= 14'h0121; // 'd289
      10'd692  : out_data_ref <= 14'h03b1; // 'd945
      10'd693  : out_data_ref <= 14'h045b; // 'd1115
      10'd694  : out_data_ref <= 14'h054b; // 'd1355
      10'd695  : out_data_ref <= 14'h0331; // 'd817
      10'd696  : out_data_ref <= 14'h07c1; // 'd1985
      10'd697  : out_data_ref <= 14'h0599; // 'd1433
      10'd698  : out_data_ref <= 14'h07f3; // 'd2035
      10'd699  : out_data_ref <= 14'h06d0; // 'd1744
      10'd700  : out_data_ref <= 14'h00e3; // 'd227
      10'd701  : out_data_ref <= 14'h03ea; // 'd1002
      10'd702  : out_data_ref <= 14'h05b1; // 'd1457
      10'd703  : out_data_ref <= 14'h070d; // 'd1805
      10'd704  : out_data_ref <= 14'h07ea; // 'd2026
      10'd705  : out_data_ref <= 14'h06d0; // 'd1744
      10'd706  : out_data_ref <= 14'h0103; // 'd259
      10'd707  : out_data_ref <= 14'h06da; // 'd1754
      10'd708  : out_data_ref <= 14'h0723; // 'd1827
      10'd709  : out_data_ref <= 14'h05a6; // 'd1446
      10'd710  : out_data_ref <= 14'h0415; // 'd1045
      10'd711  : out_data_ref <= 14'h0454; // 'd1108
      10'd712  : out_data_ref <= 14'h0720; // 'd1824
      10'd713  : out_data_ref <= 14'h03cd; // 'd973
      10'd714  : out_data_ref <= 14'h05ea; // 'd1514
      10'd715  : out_data_ref <= 14'h034f; // 'd847
      10'd716  : out_data_ref <= 14'h0048; // 'd72
      10'd717  : out_data_ref <= 14'h0423; // 'd1059
      10'd718  : out_data_ref <= 14'h0574; // 'd1396
      10'd719  : out_data_ref <= 14'h0197; // 'd407
      10'd720  : out_data_ref <= 14'h07d7; // 'd2007
      10'd721  : out_data_ref <= 14'h0465; // 'd1125
      10'd722  : out_data_ref <= 14'h0260; // 'd608
      10'd723  : out_data_ref <= 14'h05b2; // 'd1458
      10'd724  : out_data_ref <= 14'h00ac; // 'd172
      10'd725  : out_data_ref <= 14'h0556; // 'd1366
      10'd726  : out_data_ref <= 14'h042e; // 'd1070
      10'd727  : out_data_ref <= 14'h01c8; // 'd456
      10'd728  : out_data_ref <= 14'h0630; // 'd1584
      10'd729  : out_data_ref <= 14'h03df; // 'd991
      10'd730  : out_data_ref <= 14'h081e; // 'd2078
      10'd731  : out_data_ref <= 14'h0020; // 'd32
      10'd732  : out_data_ref <= 14'h05ca; // 'd1482
      10'd733  : out_data_ref <= 14'h0220; // 'd544
      10'd734  : out_data_ref <= 14'h0286; // 'd646
      10'd735  : out_data_ref <= 14'h02a8; // 'd680
      10'd736  : out_data_ref <= 14'h01ac; // 'd428
      10'd737  : out_data_ref <= 14'h0601; // 'd1537
      10'd738  : out_data_ref <= 14'h0683; // 'd1667
      10'd739  : out_data_ref <= 14'h02a4; // 'd676
      10'd740  : out_data_ref <= 14'h00f5; // 'd245
      10'd741  : out_data_ref <= 14'h062a; // 'd1578
      10'd742  : out_data_ref <= 14'h02fe; // 'd766
      10'd743  : out_data_ref <= 14'h00b6; // 'd182
      10'd744  : out_data_ref <= 14'h053e; // 'd1342
      10'd745  : out_data_ref <= 14'h033f; // 'd831
      10'd746  : out_data_ref <= 14'h039d; // 'd925
      10'd747  : out_data_ref <= 14'h05f7; // 'd1527
      10'd748  : out_data_ref <= 14'h062c; // 'd1580
      10'd749  : out_data_ref <= 14'h02a8; // 'd680
      10'd750  : out_data_ref <= 14'h021d; // 'd541
      10'd751  : out_data_ref <= 14'h06b7; // 'd1719
      10'd752  : out_data_ref <= 14'h04eb; // 'd1259
      10'd753  : out_data_ref <= 14'h00c5; // 'd197
      10'd754  : out_data_ref <= 14'h0095; // 'd149
      10'd755  : out_data_ref <= 14'h0045; // 'd69
      10'd756  : out_data_ref <= 14'h03ba; // 'd954
      10'd757  : out_data_ref <= 14'h06e9; // 'd1769
      10'd758  : out_data_ref <= 14'h04fa; // 'd1274
      10'd759  : out_data_ref <= 14'h0356; // 'd854
      10'd760  : out_data_ref <= 14'h07cc; // 'd1996
      10'd761  : out_data_ref <= 14'h071b; // 'd1819
      10'd762  : out_data_ref <= 14'h00ad; // 'd173
      10'd763  : out_data_ref <= 14'h0563; // 'd1379
      10'd764  : out_data_ref <= 14'h01f7; // 'd503
      10'd765  : out_data_ref <= 14'h0063; // 'd99
      10'd766  : out_data_ref <= 14'h0517; // 'd1303
      10'd767  : out_data_ref <= 14'h025f; // 'd607
      10'd768  : out_data_ref <= 14'h0138; // 'd312
      10'd769  : out_data_ref <= 14'h01b4; // 'd436
      10'd770  : out_data_ref <= 14'h0780; // 'd1920
      10'd771  : out_data_ref <= 14'h0756; // 'd1878
      10'd772  : out_data_ref <= 14'h0409; // 'd1033
      10'd773  : out_data_ref <= 14'h01df; // 'd479
      10'd774  : out_data_ref <= 14'h06ee; // 'd1774
      10'd775  : out_data_ref <= 14'h05d8; // 'd1496
      10'd776  : out_data_ref <= 14'h034a; // 'd842
      10'd777  : out_data_ref <= 14'h0733; // 'd1843
      10'd778  : out_data_ref <= 14'h04bb; // 'd1211
      10'd779  : out_data_ref <= 14'h00c3; // 'd195
      10'd780  : out_data_ref <= 14'h0106; // 'd262
      10'd781  : out_data_ref <= 14'h061f; // 'd1567
      10'd782  : out_data_ref <= 14'h0043; // 'd67
      10'd783  : out_data_ref <= 14'h0235; // 'd565
      10'd784  : out_data_ref <= 14'h00f3; // 'd243
      10'd785  : out_data_ref <= 14'h0697; // 'd1687
      10'd786  : out_data_ref <= 14'h02ac; // 'd684
      10'd787  : out_data_ref <= 14'h0035; // 'd53
      10'd788  : out_data_ref <= 14'h02b0; // 'd688
      10'd789  : out_data_ref <= 14'h07b4; // 'd1972
      10'd790  : out_data_ref <= 14'h017a; // 'd378
      10'd791  : out_data_ref <= 14'h0777; // 'd1911
      10'd792  : out_data_ref <= 14'h0644; // 'd1604
      10'd793  : out_data_ref <= 14'h0412; // 'd1042
      10'd794  : out_data_ref <= 14'h07d5; // 'd2005
      10'd795  : out_data_ref <= 14'h012e; // 'd302
      10'd796  : out_data_ref <= 14'h0353; // 'd851
      10'd797  : out_data_ref <= 14'h00aa; // 'd170
      10'd798  : out_data_ref <= 14'h043a; // 'd1082
      10'd799  : out_data_ref <= 14'h0374; // 'd884
      10'd800  : out_data_ref <= 14'h068e; // 'd1678
      10'd801  : out_data_ref <= 14'h0765; // 'd1893
      10'd802  : out_data_ref <= 14'h03e5; // 'd997
      10'd803  : out_data_ref <= 14'h0820; // 'd2080
      10'd804  : out_data_ref <= 14'h0354; // 'd852
      10'd805  : out_data_ref <= 14'h062a; // 'd1578
      10'd806  : out_data_ref <= 14'h0352; // 'd850
      10'd807  : out_data_ref <= 14'h0028; // 'd40
      10'd808  : out_data_ref <= 14'h041c; // 'd1052
      10'd809  : out_data_ref <= 14'h01ef; // 'd495
      10'd810  : out_data_ref <= 14'h03e0; // 'd992
      10'd811  : out_data_ref <= 14'h004a; // 'd74
      10'd812  : out_data_ref <= 14'h0746; // 'd1862
      10'd813  : out_data_ref <= 14'h0228; // 'd552
      10'd814  : out_data_ref <= 14'h010f; // 'd271
      10'd815  : out_data_ref <= 14'h0511; // 'd1297
      10'd816  : out_data_ref <= 14'h04bd; // 'd1213
      10'd817  : out_data_ref <= 14'h0273; // 'd627
      10'd818  : out_data_ref <= 14'h0027; // 'd39
      10'd819  : out_data_ref <= 14'h0389; // 'd905
      10'd820  : out_data_ref <= 14'h035a; // 'd858
      10'd821  : out_data_ref <= 14'h02ce; // 'd718
      10'd822  : out_data_ref <= 14'h0396; // 'd918
      10'd823  : out_data_ref <= 14'h065c; // 'd1628
      10'd824  : out_data_ref <= 14'h029e; // 'd670
      10'd825  : out_data_ref <= 14'h048c; // 'd1164
      10'd826  : out_data_ref <= 14'h02ed; // 'd749
      10'd827  : out_data_ref <= 14'h0543; // 'd1347
      10'd828  : out_data_ref <= 14'h07b1; // 'd1969
      10'd829  : out_data_ref <= 14'h0492; // 'd1170
      10'd830  : out_data_ref <= 14'h071f; // 'd1823
      10'd831  : out_data_ref <= 14'h0700; // 'd1792
      10'd832  : out_data_ref <= 14'h06e6; // 'd1766
      10'd833  : out_data_ref <= 14'h055a; // 'd1370
      10'd834  : out_data_ref <= 14'h042f; // 'd1071
      10'd835  : out_data_ref <= 14'h0319; // 'd793
      10'd836  : out_data_ref <= 14'h0094; // 'd148
      10'd837  : out_data_ref <= 14'h074e; // 'd1870
      10'd838  : out_data_ref <= 14'h050c; // 'd1292
      10'd839  : out_data_ref <= 14'h07ac; // 'd1964
      10'd840  : out_data_ref <= 14'h060d; // 'd1549
      10'd841  : out_data_ref <= 14'h013e; // 'd318
      10'd842  : out_data_ref <= 14'h055f; // 'd1375
      10'd843  : out_data_ref <= 14'h0796; // 'd1942
      10'd844  : out_data_ref <= 14'h0219; // 'd537
      10'd845  : out_data_ref <= 14'h000b; // 'd11
      10'd846  : out_data_ref <= 14'h05ff; // 'd1535
      10'd847  : out_data_ref <= 14'h013c; // 'd316
      10'd848  : out_data_ref <= 14'h0642; // 'd1602
      10'd849  : out_data_ref <= 14'h061a; // 'd1562
      10'd850  : out_data_ref <= 14'h006e; // 'd110
      10'd851  : out_data_ref <= 14'h06d7; // 'd1751
      10'd852  : out_data_ref <= 14'h02ee; // 'd750
      10'd853  : out_data_ref <= 14'h0175; // 'd373
      10'd854  : out_data_ref <= 14'h043f; // 'd1087
      10'd855  : out_data_ref <= 14'h0578; // 'd1400
      10'd856  : out_data_ref <= 14'h0359; // 'd857
      10'd857  : out_data_ref <= 14'h000e; // 'd14
      10'd858  : out_data_ref <= 14'h02fa; // 'd762
      10'd859  : out_data_ref <= 14'h0082; // 'd130
      10'd860  : out_data_ref <= 14'h0425; // 'd1061
      10'd861  : out_data_ref <= 14'h0564; // 'd1380
      10'd862  : out_data_ref <= 14'h0764; // 'd1892
      10'd863  : out_data_ref <= 14'h02b2; // 'd690
      10'd864  : out_data_ref <= 14'h07fb; // 'd2043
      10'd865  : out_data_ref <= 14'h081d; // 'd2077
      10'd866  : out_data_ref <= 14'h02e8; // 'd744
      10'd867  : out_data_ref <= 14'h001e; // 'd30
      10'd868  : out_data_ref <= 14'h0248; // 'd584
      10'd869  : out_data_ref <= 14'h0821; // 'd2081
      10'd870  : out_data_ref <= 14'h06c5; // 'd1733
      10'd871  : out_data_ref <= 14'h065d; // 'd1629
      10'd872  : out_data_ref <= 14'h0544; // 'd1348
      10'd873  : out_data_ref <= 14'h0490; // 'd1168
      10'd874  : out_data_ref <= 14'h06f2; // 'd1778
      10'd875  : out_data_ref <= 14'h017a; // 'd378
      10'd876  : out_data_ref <= 14'h081d; // 'd2077
      10'd877  : out_data_ref <= 14'h0736; // 'd1846
      10'd878  : out_data_ref <= 14'h0680; // 'd1664
      10'd879  : out_data_ref <= 14'h02a9; // 'd681
      10'd880  : out_data_ref <= 14'h0090; // 'd144
      10'd881  : out_data_ref <= 14'h0104; // 'd260
      10'd882  : out_data_ref <= 14'h0090; // 'd144
      10'd883  : out_data_ref <= 14'h0386; // 'd902
      10'd884  : out_data_ref <= 14'h0113; // 'd275
      10'd885  : out_data_ref <= 14'h0610; // 'd1552
      10'd886  : out_data_ref <= 14'h035e; // 'd862
      10'd887  : out_data_ref <= 14'h0388; // 'd904
      10'd888  : out_data_ref <= 14'h03e8; // 'd1000
      10'd889  : out_data_ref <= 14'h081d; // 'd2077
      10'd890  : out_data_ref <= 14'h040b; // 'd1035
      10'd891  : out_data_ref <= 14'h0367; // 'd871
      10'd892  : out_data_ref <= 14'h03d6; // 'd982
      10'd893  : out_data_ref <= 14'h0796; // 'd1942
      10'd894  : out_data_ref <= 14'h0473; // 'd1139
      10'd895  : out_data_ref <= 14'h01ae; // 'd430
      10'd896  : out_data_ref <= 14'h0635; // 'd1589
      10'd897  : out_data_ref <= 14'h05e6; // 'd1510
      10'd898  : out_data_ref <= 14'h0759; // 'd1881
      10'd899  : out_data_ref <= 14'h0191; // 'd401
      10'd900  : out_data_ref <= 14'h0446; // 'd1094
      10'd901  : out_data_ref <= 14'h0236; // 'd566
      10'd902  : out_data_ref <= 14'h07d4; // 'd2004
      10'd903  : out_data_ref <= 14'h0274; // 'd628
      10'd904  : out_data_ref <= 14'h03b0; // 'd944
      10'd905  : out_data_ref <= 14'h0632; // 'd1586
      10'd906  : out_data_ref <= 14'h058b; // 'd1419
      10'd907  : out_data_ref <= 14'h0787; // 'd1927
      10'd908  : out_data_ref <= 14'h0638; // 'd1592
      10'd909  : out_data_ref <= 14'h048e; // 'd1166
      10'd910  : out_data_ref <= 14'h04eb; // 'd1259
      10'd911  : out_data_ref <= 14'h02f9; // 'd761
      10'd912  : out_data_ref <= 14'h06e7; // 'd1767
      10'd913  : out_data_ref <= 14'h0271; // 'd625
      10'd914  : out_data_ref <= 14'h0833; // 'd2099
      10'd915  : out_data_ref <= 14'h02eb; // 'd747
      10'd916  : out_data_ref <= 14'h0312; // 'd786
      10'd917  : out_data_ref <= 14'h0167; // 'd359
      10'd918  : out_data_ref <= 14'h069b; // 'd1691
      10'd919  : out_data_ref <= 14'h0498; // 'd1176
      10'd920  : out_data_ref <= 14'h029f; // 'd671
      10'd921  : out_data_ref <= 14'h0209; // 'd521
      10'd922  : out_data_ref <= 14'h06ef; // 'd1775
      10'd923  : out_data_ref <= 14'h01cd; // 'd461
      10'd924  : out_data_ref <= 14'h054f; // 'd1359
      10'd925  : out_data_ref <= 14'h06e6; // 'd1766
      10'd926  : out_data_ref <= 14'h006c; // 'd108
      10'd927  : out_data_ref <= 14'h0734; // 'd1844
      10'd928  : out_data_ref <= 14'h0065; // 'd101
      10'd929  : out_data_ref <= 14'h0265; // 'd613
      10'd930  : out_data_ref <= 14'h0745; // 'd1861
      10'd931  : out_data_ref <= 14'h004c; // 'd76
      10'd932  : out_data_ref <= 14'h0801; // 'd2049
      10'd933  : out_data_ref <= 14'h03c9; // 'd969
      10'd934  : out_data_ref <= 14'h01cc; // 'd460
      10'd935  : out_data_ref <= 14'h02e7; // 'd743
      10'd936  : out_data_ref <= 14'h0603; // 'd1539
      10'd937  : out_data_ref <= 14'h0544; // 'd1348
      10'd938  : out_data_ref <= 14'h00ed; // 'd237
      10'd939  : out_data_ref <= 14'h00a4; // 'd164
      10'd940  : out_data_ref <= 14'h01ef; // 'd495
      10'd941  : out_data_ref <= 14'h0507; // 'd1287
      10'd942  : out_data_ref <= 14'h0112; // 'd274
      10'd943  : out_data_ref <= 14'h0344; // 'd836
      10'd944  : out_data_ref <= 14'h0755; // 'd1877
      10'd945  : out_data_ref <= 14'h0794; // 'd1940
      10'd946  : out_data_ref <= 14'h02b2; // 'd690
      10'd947  : out_data_ref <= 14'h06ed; // 'd1773
      10'd948  : out_data_ref <= 14'h0605; // 'd1541
      10'd949  : out_data_ref <= 14'h0561; // 'd1377
      10'd950  : out_data_ref <= 14'h002a; // 'd42
      10'd951  : out_data_ref <= 14'h03a4; // 'd932
      10'd952  : out_data_ref <= 14'h0291; // 'd657
      default: out_data_ref <= 14'h0;
    endcase
  end

endmodule
